BZh91AY&SY^j�8�9_�pp���s� ����az�              }               �      �     
     DB��  ( �  �       @j�Q�( ���(4��Y�D@�2;�3�þ���}�шuI� ��A��=�8 �ťR*ɠ(�8 �`�.CEQYh(��RF@]� � Ub� �Z��2�S&�J  8JD��T�vҀ
�0 8 �-IJ2���$gn���.�B�Ԁ��@�
� һ� �۩��  �d$b c� t�����F�]� �p�T��h�n���RXƊ �AJ(�����@�@��*� oW��{��Ƕ� �n�Èwe���u����x z��年\m8 n,��2�z���J�h����%wn�k�n���Vv���-Hť\  �PBP��(�Y�@=�w9�s�����F���}�>__y�oI�׋NM�1��x �����ɥX�� 7��r�ܚS�R���(�g��&�[�.�x�y�U���)��>�]��v�M���ͽ��u� ��A@
UR� *w�����NYu��ί;�^�� 7}}[\��N�c�+��z�� ���O__}�_  f����m{}�
)�J��|y�x��N{�kۼl��@S��Ժ㻫.,|��;�W��    )�ShҩT�4��4��������UJ�� 	�    "x�T�F       ��U*U h�h 1   i�d��J�F       D�R�2h&L�m=M@�j�d�(�=O"~�������������u߮�����%  �2��� Z� ?�@ ?��� R@?�@@ '���  ?�/���� g�]� ��O�@��I���`��� �Q	�!_ۍ:�}��n[�o}������E�ծ�2u�ƪ������\
 o��K���\�
��A$/Wf��Z�v��5	fe�kp9�ZT@�˙�:A$#��T���4-�UI�I�(��m��0J�JJ�A5d�h�j�KB�P�Y���Ÿ�j#"�7Vz� ��(���ؒ	 ��+K�U�=
��E(2Y*���S�,.&B#��/Y���׫P(,�uǆMl$$aP:���?H�JJ�IʩI#�����5OC��\Z�5��7�2��.5:�nđ�l4=I"�}�s��lvdF�n�5�N�$��	"o�v@*����?@�����wY���4������%H���0�I�W�m���$*�L`�����J�N쮁PI�
������������nk[A$
�hn%&Fo2[����G�k$t�͌2撬��r-�$di!SF�r
�c#KPI�A$Z��y�vp�s�ì��wfV�K�H$�oG��A$Cu@QPM�.�
6�E���r��*-�e��$D+w|7Cq��A�eǋQ���F�E$W
��������Snh7�ɛ�;�XU�A�\���Y��Ws�H�o96��I��;��I��U���1n�\�dH,J��5/T�������np� �TZj%n��.�\kjA%����H%@�a�ۂH%U[�����h�V�tHVJ���6A.��T���$���A$KJ��V����Tho�V���`P|\C4G�l��-ũ�$�K2���A$6C�
� gsaCPI�U��@0��@(��+�Q#P�F���ɨ��G�m�S8\6B�q;Z��K�Ƣ��;{��������B��/����M�H�����굫J�v`�	"���T2�[2�n�(��j%:�g�X���-U4l�Qf��%$�8�d�^U	 ��{xm�2�	R��D�`G�F��Ƚr	;o�D��4��,�$�8bwT'`�@Ѽs���$�Q�7�TG+�J��$x���ކX|5���"Qv�BrYS|��j�Q!�D:wer9����$�TK53[gwT�B�����g	ǩ��DJ�!Q�NH&C@n�Zjh��$��TA$A%RM������:$����E�Q�Q����Ĉ����&@��D�-�Ti��!�۸$�H��H�
��3N�*w ��7��%i��Hv7-;NL�EA%pq����ե%J�m@��Z�H'e!PNj�9���$�9{���dap.	#�_/m��TE�k/*�A$�I��-4�N���EA$���Y���H$��Tp5 ٩L@�]m�0�5����8�I��4]���{�H�Z/�Ԩ�j&�e�騔^,���iT�֐ʀQPI^�w�*�X7��tr!Ubd@>����M�@aV$���#;Ĩ$���%����T�C�Y�P�(�QsR�`SP��vi�Ө�ɬ�2 Qڢ�+�I�@����	!�[�u�	UZhX��D�%��!P8N�s���&塺��y��"�	�Ą�E�3���rm�T�02��q2	#�%D*�F��X�A$o�}�E��ɴ$M�Cv6�x��H�J�\ʑ8՛΅� �J�p�P��W/%8�u��CpM��rl	ʔ��$��P�bT
:h4�;�A�L��bH$��I (�*��4�`���R�B�!����z��iPN�\/@l�2�����{�\E�y����$�|�T�te��y��:�q��aR���`r��/�P��#��h�$�v�8$�H�s7���Z��#f�/z��:IŅ@�auЖ8H������l��dB�t��PND2�h�L7����4��!�T
�����q,2�Ikmh�-В-4N۰�%A7WiIY
9���p�4o����9/n�Q\���k�æl�z����H�؇�@v��/�*;��$�m��M��m��ȝ�Q��p#����pI���v�*A9T$�r��P�/�iPICå�Ut����PS׷�\K��3'
-�� ���,�A'���Z��_��nh(7/HTk�:P\aj��Q��P�[��*k���(���x��[�� H
+���^v��p��L�H���A��6j!u�*FD�9�j���5�$Jtd+8���PID��٫��h.	�&���lf��PND2������nj��*�
�q:�^m/�A-�@�8�I)7�&r� ��obr�I Ԣ���dz��\lf�*Q$�n�I��T$�IJjO��$�H&���I�I�I�I�J�A$A$A$A$A*�I�I�I�I�I��K�j	 �	�%�$A$UBH%�$A$A5�u��=�#|�F�0�*�2\C*��N��	�y�*ovY���A$cZo�6^p�i�$���$�A5.	!f���a�n-<�N]�gCzhupI)
�� ƵsfA���i�$�s/����Xb]!U��}�c �2o��1n��a������J����N� ��W�V��$�kw�g�M��E�vI�Ѐ;�&�Ǐu������L���R.��2����\�G!�T�P��j	p��[r�T�Օ����7S�M�9� �.�aP�a
��&���!uy��D7]pypI(oFA.�I�I�I�I�I��$A$A9�I�J�U݉ �	�,��I�I�I�P�	 �	 �	"bT�A$��UU���^u
��l���`� +{5�ݩ	�k;/[��	�%�Y.&�Ts{����8
��7�tjh��I*�r�sV�Z�H]�$���0
��c���Y�3�f�p�h�����[�M�d*�Q&�N�`T�4�6Ѽؒ]�$�C��)��K�g~��9�G�R��Z{���R�q2@"D�wKt�>l��YeWM�Ph*!��ݘdB��]kqi���TB�)w|�,����MF�����flͦ*n�gu;ɾ��pI,�M6���ц�����i5�=
�������	(K�vvl��Sd�F��:���$�H'!u��� �*:a�oE`ȝJ��jҷ�p
*��rd�r	 ��H$�H$�M� �%%A$I�I�J�n	 �	 �U	 ��M�$PI�MA+��7�I4�n	 ��?=Z�H&���Iڗ��H��{ӹ(��pI���@TA$o�r�IpI�h7��x'"�j�ͅ�
�iPI�F�Rj�\ѵ�K�v�te捚L���U�\]��I�I�P�	 �	 ��H��0
�T�����Q
�_�F�+�"q24���v���IC*�l+�p�xhj��!��E�
�I5��@��v���6�}�I�I�P����*d�H$�E:�JB�P嗾��A$ij� �\�VV3��&��@(��E+T�u�Vi
�n	�7��*�$�M8�A�TD��2	 �T�-��Ʈ�h�v�WU5���J�wiFC�TM�A$��l뉱�b��*$K���]�XP\�J����/`LIaʮǙY���.	 ��7T�R�zpn	�I�9�rA$B갱��H%�%�7ۏ��c�&��)ĸr-A$����/���v\��T��D.�kQ��	y�ӗ�sF�y �Qz�"��]4�\8A$+YT@.��
��%��̚a����@*��x����p����|d�۰��Ԡ�\t0�5]��\>�D��(�gD�N�;W
t�����#��[p�\��A%����6|\�%A$�-SA	UNgJ��	7����VĐIɆ���4Ca��Hj�.˅t�G>�H$�H$�H$#�F��QT$�w�:H��\F���$�H���z��NMo���t�R[sֹ�:2	'�K�{����O���_�ߞ����� h       �8   	                              �x|                                  �޼[@� ��                              p               8  [@   l                           � �        �                ��     ��           ��  � FY�� +�.� 'Xm �� OY&���n`/M7n�Zܖ9v��1ԯn��'hકJ�]�VP����U���q�m�m��h �M~�`���-�����|���� m�      mͶ -���  �j �� p m������ �&Im�h   �e�춎8 hm.`m��  � � [A �ٵ��l�� �͖�  '��oY]�6�l&���V��� ��!pm�fS�&� &� ���mU�`  �  8        '3   ��x�m�K(�7m� ��  -� �N���Lۛ6�.� l  lm�m�  �6�  [@   t� $ � 	 �  iY#m��� 6�m �N ත��    Uc���-F���h N�� m�A����@ 6׭�lm�  qm 	�  � Km  ��ɒ '��  6�7l���   ^�[6n�[B@�6�6Z���m	i��8e�v͇6��Ĝ H��  p�  ��	 a� H   $6�'nv�nX` �$5���m  e���||  6�<�֜��ڹ  [K���� ~�}>��o��  �m��8    �  @�� h��� ���ۮ�� ����ӄ� ��  ,����a���    p-6d�  �   �K�Rк-   ��-��Yx6ۅ��    �T�PR��;s��C���S��Ʃ������^�^��=]H�́��;m�    >>��6�m�   � m�N�� 	�It  �[���yt���=*�H�CP�/�G<J�;`  7m�ض�Im�H 	����� km� m� ��u�엣  M�f�6�6�M�h  ��Ŵ a��m��  -� ��    ^�   H�   -�  �  ��   �   -��` �     ��  l p �   �@-�����H ��9���l$-����$���   v�    	���� >��&/I+���U�v�q�n�N��)8����޵'�ۃ�k�I@��c@��u_e�%�m	6�  [@   �` I0 l  Ui   a�  -�lH ����   6���`     � � [@  $ h  o� �� ݖ���e�Z�   ��h 8�k t �  �mm�hm�ٶ���	  4�hpm����n�8 ]�TP�f�h6M�e�vպK���T�`�  �  : ���  rt�E����� <���� t�\:� �	+����,n�pݶK g��8���W W]  m'V�6� ih�[F��l h6'[@6��� 6�	 m��Hݶ $   �g��J6� ӖА    v�� ������� �  � �  @� @ m�&�=� �K[l6�    �,�m�nݶl��$,-\�n<v�  �� �M� ��   ��n��� p     [@  �p�-�   �ع� 8 �vʹ� Kn� ְm�ړ�4�� � p��AmE|	���    I ����m�h�����h2-�-�l   HI&,�@6�H	I     ݷa�l �6�( t�� ��vA=$m�`N��m�` m�`,0���j@඀ m�m�I �&�� �  -���m  � �8 -���f�i2���3l :ޝ+�]7`���I�e�  ��(!$�Ԗݶ��Yv�-���  ��٦�  9�`�l� nӠ%�dݵ�6��h ��H8�@�� oIxv����l   	ۑ�sd �}��@TQT8�-�T�m�����e:I	 �6ٺ�j�` ����l����M��..�W�UT�J�ԫV5���5),�����p�2���&��W6p�M�m�l�M�8#�m�V�#m�������� �ֲT��8m��j]���Usg��-�@��L�L Y��(  x6�&����`m�� �@9�ۦ�n�  �@  �m�������U�iwe�UP�X�,�ڛ6�  nݰ-6-�hm�  $K+l@
P   l�Ͷ jl�w�ڶm�H[G�	mr�6�! �� 6η���m��-�!mp J2[m� Mlkz� h���m&�k�l[V���-�)rM�-�8 ��m��g[)�8ֽ,6�@H����kh8t���"Y@n�q$��6� �K��`Z�6� H A@� m����`  ���K.���H�l	`�     kV��4Bɖ�m ps�@�  � ��q  4�H8����f� p8  H  pK4Z�+�*�Y�v皕PF� H�۰���"tv ���������*����s3j�[ Ml�Hڦ�-��m�H���u�i�^j���wh]m\5��e�� ���2mp$ 6��ր�kkm����86��նդ�q!��M�p��f�P�  �Y*@;m��ڭa`�l �$9m�d��#m� ��    �kd�L$�  2 �������Ӟ�Ӆ���2�6z��7H�����m��� �� q�k�.5l��ց���v�]��    HڷkXd�e�5� �n�Ȗv��f�:�Ҷ� 9m�[{e�������[@   �>ն��1l�� �k�^�m�f�  p  6Aݻe�  ��{m�nݰ���l�P  ����8   p��0 l�M�� 	ky� ��@�q�Ƶ� ��ޮtd ��>>6>��XZ�U��d�@���� � � ��  ��U�`H�  m���[m�  ��="� ��   ��l�ޚ\l 9[w��m��u�浇  �6��"L ��hl��UQ�6���. ޼�h �d�dͰ #Ep�ݶ���j��`0�s(].��GZm�  �I@ [�� �����m�#]�l�]6� ж��k����  �l� oPղP�   [Nm&��m��� [\  K/  M��[��"P8� m� -�w�� �z��  [@ ��  -� �@�@ 8  YTz�kX         �I� ����    h �  �dp[@-�� ���h�  9�k�U6�x�`  	e     C��< t
�P���m� �K(�f�l�> �,�j
��4�Ͱph����w{�����U � {݉���������D����Q�)�e���O���@
lQ~�8��Pt�A��� 'P�������i�c� q�� �i�qx*/l,��(�U��0�UbB- ���XD�L �	�# $E�A�D$EC�����J]Ѝ�GC��"�b�X��T��B�LQáh0Q"t��AT!�bn�ϕ8�|���V"�*����\8���z:Q ��A�S��X�F��P�dU�Q4T>�K@Ĥ -CAM}�>A�pj�b��� [9��}�A31$B
� D�$H�E�QB	j��~~KD��>Ҁu���E�]� ���,� H�mU��V��P-���1ãgQ6�ڥ
�b,�2
 D���)ФJ~Co� `$���Z���x�H)N�=Pv(��(i� pKڀl�����#"������V ��C�b||�a�BB����N/�&"Z�@u�)�@>� ���@�/���   �^���7�W�_�������hD?��u!p2�P��Dn
"A��B�"!LG�{��������� <H$     m�     ^�ְ     [@  ��      l 8	  �`6�� WU�����ĝ�n��I�h�J�v VUVV�R.)�݁�m�7�5�R��yѰk�4�'[r�V�Tځ�qӳm1�{mmP!�ڧ��ٗiy��H&�ڴ�*�.խmʉ��v%�6��<	�:�$-���l�y�At&�uյ�V=m�,������&K,�Np��5�m��l�) T�m��ѧmD��NuUu��w-��- �ԫԩ��ʷ�n��Ͷ��	=BN�]�[6�b8K�T�X�֤-��ְ�`-����n[���c���z�ۭ�N�U�vN	��M���YUWTTdviV��.e�8���M������IS&��R�Q<v봝C�ON����v(
W�*�����vͧ����K�ʠi�N�wk��)$��V���́�յA<u Y�nKZ��\��\��"cS��R�ufwP�Kz �r�����8�Kz@�c��T�3:����gRlT�<P�vE����ںyZ�!��Ć����i+a-r�v��z�5Qb]�\fu���h�r�bjګ�rF�Z�wj���J�;���k�^ݻ�q���T��<\��k6���#�dP��a���i�]kv��\�&��&��C�tR�U��:��`8yR9��(2�y#�avVwe�xs�v��λq��S�����6���ʡJ�ɰ�i"�������ٕ�vri8��G!5��.�B���p�0E��藷K��lkx���6�J��V����vP�`��J�ɶ���X�ݗI�m;������H񝔚�}��7Y=�<;����U���L�U�i\񋢶�2 J� ��J�F�` �^�r��
��F��UUS� Ւ]U7wy�EVwu�^ )�?��� �!i/D'lE����D�]#AdmD1@�-A�6RZ'UQ�!�]r^�3l��Slm�m����yfmg�V"��
v����� �vV�a����m�=s�f�&���\X�ݘ��v7z��hÜ��7I��]⪗��I9
u�5�.��������v�]�0�<������`�D9�:k���j����ۅM$m�!�i�<����T�isּ:'0����H�����r
��E�MIu*����uuS�yP�vˇ{yv91�p����c��87'n{o�0�����=����Ӿ�dqos�]�s£-�m���P��|8G���>���;�x��%Y��a���6([�������dqos�\��(b��#�p���bh$�H�g����C~�	���ŧ�p��ӌ���`��bl�����P��y�c�s���C�q��L����A ����D��h'l��;�%�g��4�6.�v5�耼��9ݢ�Т4��\~��߽������5k���10g�	L�����7���ffM#�C=���8���&~��߿8���Ȅ���Kg	Ldqos�\��(b���1�9��z.�r���P�^�m��?{����{]�w"��}FG��{�2��%��a-��i��e��3�>�Lq
���>�=��p�/��[~��vN����)��Zn��{c��!��8�������\��rN\j�b�o"�O{�G�9���{�a�����@�L�#A�I3=��g������.�KW.���{�,���8�O!���x���q�~̈r���C�q��h�8x�a�L0q ���.�KW.Ž����w�1|�`�)�AlHq�C��g����_��8���"�?~�����M�x0�����6�:<#u�E�cWL��ccZ�坫����j���$�� �Yx ���c\_[<!���x���q�!��3�q��($1����i��/�2�]�w"�|��8��xK�]ί
Ж����0���8�?��D9��/�1Ÿ@�=ȼ	J�V�����o_.��������V��)�����C�b�X�, Y4"%+  � @Z��Z�B�H!��Z&�W�z���}�@\O	L�fz!ϸ�E�q�.?t��Z�p�$Gܐ� mX\q�kv��g��4^[�s����2�qq�OA�
��ቲ��r������c�s���C�q��q���0��K	#l�|�dQ-\�G���ժ���10p�vK�N� �#�s���S��ս}�`@RA	�z��W3������_,��#�-�LG���(��w�1i��#�3�3}���X"�J(a/A6��_�⿳��w5j_*�����=||yP�T�_�I$�I%KU*��+U@R��4q�e:n;N�nq�vm��-�`�.�ot�H2է{#ڤ��v�y���g��	�mr�C����W�v���Pn�(�2#����Ƀ�crrq������">9���u<�#b��g�͌��՝ϧn-��9��	F��9֝ڞ��q<�mج�޷;�Ӟ0EV��Gq�z�Q��u��N�(�Ʈ`Ȱ�w����)��f1�n�8_&�Ru���m�C@g{]���pڇo(,�V5���%���������./�1�9��z/���_}��_�@�(��ŀ���6?S6������*�l��}�B%��$���zYn��;2侸��2z/�����]��%���8���~E�!y�i������,:b����./�1�;�=��p�a��0��O#��]2(��\#�~��]����~�����]�'�C<s����I��l���l彮�zu�2� D���h9�Ƹ�Z�-��$bz./�1�;�=��]��E���Ah��<�̴�qo�}|+��B
����_/�����UJ�k�S�*Gz�@�̼	c�-��_�dqw˦E�˄qo��"���xT	`O�Pd4��*~�F�U/��!�t����"�p��{�xR���-'�D�\�G���(��w�1��'�w��c6�m�t�;�N�z��9mD�ͬ-�V0�j��CcŝƜݮ���spc�똣�~�t����"��]2(�˗�ӝ��@2Y_�&�LE}��!�{��\_�c��~f���E�>`f���K	#	Xn�W~ټ��o��o6��@,����"����A>]�GE�)�踿���d�_r�E��K圹�MĶPI1[�����0�7�p�����qqɆ
!xX
���q�}�6�F�z�;;����vS�����r���� ��V0V!��-�����"���28�˗�ߗ�E�Ĳ�,%�-< ��1o��~Z�U�^�z̞��>��j����xY��[��4l��p��cs�꺰��꺱�"��D����a���!�t����"���280����ϗ���=�p�[)/�I�1w��b߽�0����8�}�'��_�������9��݉��c=t�k�E]�X��Xiس�s:sZuc\mqŵ�]�(a)�Qq��Gǽ�#�~�3�ٟ�k���-hq��M�h�1�M�����C���}˦E��8�hgv2KI���%�)1�ſs�]����@$@#�E��)!�?~�rtj������
c�+0�ef��ĄV0�1$}�{��*~����p��ߗL�+��2�_aZx$�A��gN��z�����C��f���������IQL��P$`��D�"�@�"��ӣ����  � 	:�j�	� �τ�tn�y�5͑{���n���:�C[Gm�T.#B&�\llۮz�pCӰۜև�ݸ�;��v�s�.7;[cm���mۮv'N^�sW(��5��х�mu���܈rj��s۱k\s��g�n�m�O�pn�gM�.�-�`ێn�鶹{G�����
�Y+9խ�v�l�[���YCu=�PN^��6`o�{�y��I
.&;�Q;�#��Y7�g�2	�htuM�C�i��F�V���nyl8��؏W�28���"���x����(�}�@v'�����2َ!�t��[�lmg�l���l���G�y���L�@2��m6�(�z�����(�?��D;�=�����8�F�G|��(�=�[��K�3?~�zXt�����/iq�)��?��D;�=Ǻdqw��"����֒Sa��z���벍���7�;�[b�.e�v�0O:�^G��b�) �D'��Sg	Lf�_r�"���x�߽�����5���躅VB��e«*eʫ�z����f�>���^y�"�Z�Y[���k�֒�Ȱ��$��S0�>�Q=���wL��}�2z-��p<,���xQ)�����ſ.�Z��(b��OE�1$�fDJjz!��'��L���{�|G�5���<~,��㒥�'^4�1�l	�a�%p���3q�!�1�K�2u�D��Cl�K�Ɗy_}��!�{��Awr��wt����8xbe�,4VS��ur�Z��VG��E��|b�Z����d��'1=]ܧ���k�OـpИ�C��!M�)�2%f��c�/bo9�`��h[B��I�Lb��12�R3Z��Z�	�J7�i�2�sb�
V��F Bѵ��H�[b�K]R��m�P��,�zB�ir��k���h��q��-��)eC4BT9����((�f��ۉ�f)�]�)Ǔ\�/,�U�@�xCC�.�(SaH�W>>P(��h6�p|>R�v �����O.���T]4�^�a���*Z&��� t��B�V��ƏGp������y��_�����.�7.2�	E��\��� 
�����a�d{������r9@�W~ߦ�Cp9��{޽��t�-g���mB�-���c���.�A+�oV.��tJ��+��]*=�ŋ�\J��f�b]+��^����V�ٔ��s�rq�z{=�ܕ��c���w�v�{V;Otv7�sK�W�Ȯ�Z>�Ψ.�A|��y]	tP����tK��Y
���#�H�#�jk�p������uv�M1��ڍ���(%�B��lX�*�T�7��]��m��r�����V�DM��2>,�˓�)ah�E���\J��ݝ�.#����9O�{C߳�M=�G�B�~��et��A|�ޱa-K����(WJI(V�3oJ�t�+�=����y�g������/�>U*�!RDZ�V'�F�U0�"��:Q	�{;${Ǒ���Ң2�Zm]���ҸWJ������P��&, A�}�yC����g�jG���V�i\)��x= )��w-G2�,.Dsn�{\��\�j�v��k��L^E��bUUJمُ�E�v�Cr�º(U��y]+��PW���WEºT+}�l� $�B�#Q�u���i�p��ƽvH!�+r]�#Y]+��P_l��WJ�WJ�n�6�t�.�A_����]*��]\J���Z�d-�+�de��B]
蠖�z��]D���6etPItP���.�p]*�ՉtP��	o��֮8�rAܗ��At_��?s^W���E
���磐7? �;B�~�� v�!������D�����"�E��ۓ+��]*=�ŋ�\J�}�z�.��A-�f�.��((��̮��]���ڲ��I	!�EH�X!D�"1��wN�����?~����  7U`�Sl6ٲ�Y�I,�n�;g��s��`s������9�n/Y)ַ*r��L�4�ɜ�' a"�z�)�ݘ{`q��Y���j���m��t6���6r� ]�[�p��]����77f�����H�(�Kq��'K��T�����x`�\�ug�7��<��wg��S��{v5�l�m�U��{q��d�ֵ�V�[<�Km��UR-�� K� \̴C36w\흛�͹9+�I��a��[�i٧8����	ۻ�w��-]��^�T��ӨK��]����Ұ]���ي�(%�B��رtK��P^�e�81;��n���.��A-�3oJ��.�AG��et\�W7u��Ҡ�ws�?��b)�����(��l��%d�n��X�V�PSg��A.�6nᣐ5 9�}���2<�@����.��(/�z�6仲K���ܚy��Q#Y�z�r���+��p��n<�@���9C�S!�g��z,�^�/-$n\L��J�r,]P�r�{�����_}�z�r9@�e��f�Cp9�g������|V�:�~���D�pdK��{��[�^q��U�{/�\�V��u��}��:��=����b�WE�=�Ջ�`�%=7fWE�]*l݋�I	/��/��{��ՉtP��	j���nID˅�r^.��((��̮�*���K��`ԋ�e�1����C������Ҡ�wgP�Eº(%��Ջ����(/&�Lpv��etX%�B��y.�1t�/�oV%�@�D�{����գ��9!��~�]�(W�I~Qs�~QKE�%����ó�CP�߿gH���A/�ub�X.�AOMٕ�`�D�(T��"��&.��0^S������r�jG$X�tPJn�鋥AtJ
}=��=�p;F���^�@�9�~��8@�WE�ۡ���$���j;Wn��=��X����x�th��i:��0��b�=�{�gv��嶮�E��t�D������K����{��4v���>���i�;�J{��J���K��U�E���wnL���(U���]B�T����WE���b�X.�AOMٕҰK��G�^�$�Jܗn�kD�.����ĺ(WE���1t�|��Y $��;P�g��<��]*��^.�p]*�Mk�����ȣ.�b�WET���ެ]+�()�2�,�W=��.�p]����ĺ,+��^�\j��m�8!7$�Ҡ�%�ٕ�pK��%s}�D�.�{�:��.�A-{�X�V�rs~���G��m3��"#(C�f��ϖnˮ�uy*cn���&�����C}�Ʈ���YnL���(Tg�^.�p]+!���h9G�����h� �u�`��l��%�B����v���ը�j�G��\J��ݝB]*�WE���b�X.�AOMٕ�`�E
�����W�U�|Vy�~�&��B�qb]�A)���.��((��̮����F��z�r���+��p��n=�V�C�ˈ�Gn��X�V�UUAOMٕ�`�E
�����.�Av��CQ�8�X�E�-2 ���H�`@߽�f��!���Wr]�q�ܒ\�+���E
��׋�\J�W���K��]׻Ջ�`�%=7fWE�]+�f����	��d�����j[���o4��wv
�v:	�ʜ�eD[���(Hܸ�q�ǋ�\J����b]�A)�f�]*�PW�{o+���E
��׋�\J��{����."ژXf9�K��]�f�b�P]��H��ߦW��/�
���x�%�t�/��V%�e"�(%�ۍ��@l�v�$�Ҡ�%g��.	tP���x�%�t�+���%�p��	}�z�t�.�Ay0�58�c��m��+��.�+XVC�ǋ�\J����b]�A)�f�]*�~�),�7��|.	tP�ɬ�&�B�hR;�.�r�B��g���d {���C�()�2�,�Q�{^.�p]*��{��t��/� ��m�/2�UWR�s�������1fH��x�.��w.๽�U��ΰ^O��g�F�:�F�y��$mY�E�󗴎�R��ݓ�0e�z��.6wHb霻vwknv��`z�!a��q�5ّ��9����X;v���\��K�{n���iܜQ�Q�ȵu���݇q�0��q���ə��u��-h��1����vbʶ9%���/�t��������*=�[qۣ6ݮ��C��|�֞wg���9.�8E-���+O%�`E��Y���h;G�����~���4vT�PW��ו�pK��\�k����E�X+���c�WE��p,F_�5-6��ݸ�t�.�AOMٕҫ�(Tg�׋�\J����b]�A)�f�]*��PW�zް��;��!�y]�(U���]�T�n��*]�f�b�P]����+��.�Ǟ���J�%�v����ĒU���ĺ,+��S�͘�TD���}���v�؈��g�~���r9߳�]�[LWdQ��%�p��	}�xh�r��� ��=���j!���{oD�.����ĺ,+��^�^�"�ړ��ֻ�i�N�dϹۆ�3�@���[�
s��5�\�}��{�㧏��nrL]*�PW�{o+���E
��ׇ n�B��{W��A;G���O�X�TD�����"�qIe��ۓ4���dr�_z�r�@�!��2��K�º(%=�ً�AtJ
��m�tIpK��{Iw�ۻ�V�%��.�p]*
�7q�t\+��_lެ]*	R���&WDĺ(T_��tK��P^�#6���pCujŉtXWJU���1t�.�A_����]*��^.�p]U�{��b�/�|,�j���ˈ�Gm1��t�.�AM���+���ET2�_z�r���;~�5#�a]*=�ً�B�TIRU鷽��!e�K4��c�\�����Cjy7^��;�ֻ�Ƥ�wO_�wwk�q+@��N�^W
�]*��^WJ�T�n�et7��u�g� ;�#��~����ܮ��Aj�F��+�D�ۗ�Ҹ.����tU�t�T��f.�
�PW�{o+�p��s}�+�%�t�-g��jڅ�[S��2�.ҡ_lެ]*#�Ͻ��F��l-Z��w�oժ���Ay�{�]ҡZ���nIR��˴9&.�Ғ����y]�(5��ף�7G!^׳�O均#�a��IpK߹�����Ɇ��q4�n�NG&WDĺ(T_��tK��P����{���5G#�Ͻ�9G��Wu��O#���}��]��L²�&G2��;E�a�hyM]��Orc�9�܁7mO4r<�[���$�X�Q
�H��y_�E�X+������WJ�{��Ջ�AtJٻǊ��b]*?��x�%�t�/��z�5.]I$�谮�	O��b�I+�rB���Zy��25�}����#��k���Tq�2OnJ��{%�i�wn�ŋ�AtJٻǕ�1.�G/���G n"�r9߽�A�j<�	O��b�X.�A\���z�Ewq�e�V�Cp9���o^�����#��ڿ߮Ð�y��g�h�r� .�j��{�ߞWDĺ(T~/v9;�[�U�U�h�Ñ�}~�!��_�{^.��������/�_
ǻ�b�K��P_�s��H!�����&�����6=n�ۨ{F�n�c4s����d��w���Yn5�K�l��^9���p��	}�z�t�.�A{7x�&%�B�����UU�=��v:�����5C }�����Q�1t��PW�{o+�UR��E
�Ok��,J���ަ���d��ᣑ@.���ޕ�LW.&;���<���tP���m��Ñ�v��CQD^C e��f�Gb������\+��n����w���WJ�t�UIA^��XWEºT�}�p���y����zy�!�` 謞��y_�t�-�F~��i�n��tXWJ�O��b�XWJ����y]+�tP�d������PV{��et\+�A�����q�h,�,kB�Ȅ�"��K7��(F ��!k��b:A�ќ�������B�5E Q]XȰ��I�'P�P�=%�w�1Aȉ��t0"���m!��p�1��p�(��(㎐��H��+���k����7����k�lMt�M�h�
V�(l�����퀅<�w�$����V�6	"F�aJ7XH<�WQ�o*	"KN�)�c� R��*jb�Rh�<#bc����$K�-�D0`���VA$"�$@�{����w�;ߞ���?P I#�           �|���      [@  ��        @  8m��� �8�t�-v��p�'�-uɨ��ۇ+���`�6����b8��v�q�^�o[����g`���V� �.�F�)mv�fׯ	5��6�a���sF�΄ؚ�N�p7ga��#c�UJC�����32�Z��	Ci�H�e�^�Cn�z�����$;��;�������9\ݠvZ�Wf���t�X�Nj���涞�md�J��U�q​��&uC�$�w)F�f�!�^c`����NP�b�p	Ԏ	-� j�Tʴi��� ���N��۔v���g�s�����J�PS�.�gm���rG S��Ҳ�9Z�f���������+=��R�YC#�Z�Cs�K�ڮ'l1�52�Tjc8�檎�ހz�V��S�� ୪�g�K��Z�r�v�ېօ-�N�jR��ɘbL�WWm�����e��j�� ֦��O[�G7U�`�V}{:Y�"ޱ)y:�z�D�i�`�/i�	��۵S�^��	=��:w��hgn�[�[3m�b�1{Tp�����NE�J;}wͶ�n�n���m��M�����ݞ�k�6� �5�r�HmJ�fU���#ܖ+lj:�0��b�^n����p(Zn�5��$�p&�8jA�������[mJ�5\����=��A��X�K��y���0Б�DO;T^^�u��+����k�I��:�\�S�J�ث*���vֺ:�UV���{O (!U��WJ����U�Bi݇8)ǳ���B��;anY]��)@�@l.	jU�H[�
�eS��J�p$�% lQEʧ\n��8.57J�QE��:%USa�:%��V죵Ta�������T�N����U�����/��¹L�ee��eY�GI��Ώ�C�pK�4D�� �x�m����f�M�T�u_w���{��ӽ��qI�  0 ����ݖޭ�u��_��g�y���c��`�<���!�۵!�G*�nû)��g�0����`�Ϟ�e-�3��>R\e�6n6��Vj��6�m��nn�pn4g�p{s֭���r����;��*�{�7�]�8��^h��[�p��qיM�N�v.�[��v��xss�i���v�۰k�]������/<���.ش��<�p��n�@q�Hm��g�]ڸ�`��G�ؽӃ�;����8�����N܇�ҡ_���o�<����Q�����\J����b]�A)���]+�(/��U�ܖ�#��cr�.	tP�g�^.�At�+=�i�WE��昺TD��=�y]tL�H-�FԹDD.Q-��X.����K�º*?l�°T�߳�y]tL�Of�T�����hk��VژXcɍ.��tU��i��AS���&S~�m��*TAz~���XWE_���RK�E�����¸*b�����&W��oCp�n�}��9ǐ���>�o�� ���r��+*��'rTQݒ��(W��z���nb��TT6J�/5��t��\ܹ�n�RGWE])�_��V�1|�wA�j<�u߽�7��s��է�y���&�*Z��<T����kG$�"�"�m(�EZj�h�BQ�%N���j���h�r��ו�WD�o��U��L]OM����r�jI$ĺ,+�����\+N��i�N
)$.?g���n�¾�{Z]
�帬���Kl�n�C
��/M�����&S~�m�
b������y�!>�~����;�����`��j)����&W��^*b�LW�����p�����1p��+U��<��]*T�߭������S{V�=�l�{�9�l���e�TmRc����:�0�F�V�#nܾ*�t�.��ĺ,+�����\+L]�=���WD���k�L\)���kr�4���+�1��p�����1p�*b��k���R��|(S{{��V�1}���K��tU���^�.۸��rI��`����m�tU�2�=��U͏�'D�BTP�Bh��X�o;ƗEº*��i��AS��^� �r�s+�����߶�V�1w�w�]?�6b�P�j�.��+���I���N��.8�S)X�>��.�$�j��b�T1~���WE])��m�
b�z�n�8;%��;����C��ĸ��n�e�g�oV�noI����Fe7M�;t(��ĺ(WEO�M��T�p��o�O ���z�~U`d9����it\+���U������v�܆.L[���]tL������\)��Ͻ��2<�}�=�7������ ��Q
�LP��I������j��l�7r�p�諢e~��^*b�LW��u��p����b�PTž��WE]+d�F�"�+�q1˒�:��,%�>��������h�rß}�M<��hC몍GMi���^*b�L^^��hk��6)��d�it\+��y昸~T�HX*�]B/?{L�
�&U���x����ĺ(WE^Z��j�w�D�K�v'��uoAr�cgYΞ�J�Ca6�&�th��G���\'^�c�&.L^���+������׊���{����D'a���z�4n9���+k���'m�mɕ�WDʷ���:��p�״�ǐo�g�F㟑(r-����ej��0��*Z��<T��|���Eº*��i��AS߽�+����o}zb�
b�?�����d�&%�2�*zl� ���{�etU�2�=��S
b���D�.�W�w����Q�Վ�1p�*b{��4�!s���}^�C��}���C#�7߳٣q�7Б"0��\ �P�9�P� -����{����w��o�Yo� UeR��R�U*��㠙����6A[���M�81��$�N�G��j�L�Tr�:ӹ��KPn;��l�Mʣ�]�0���������'�ݻj$��vgB�tZ�,`�;4,8�tDf�ۮ������)p!X��B���nkG.�뵼�4[Z�Z����F�4	�����l��]f�auO���n����a�]��sY��m���mUUUKa�A ��뎼fp�\�l���\���e۴�t=�n
8�B�1H�N�C������
�+���^���+��=��y�^�:)ʬA=��etU�2������\I�D���`�S���K�etT��ً�I� ��{�s���<����~��*
b�I�w.�2�q��%�p����צ�� �/���O��=�F����\)�߷?b]+��/�������
ܓ
��/}�i��WD��ٛx���1^��]
�|�L\*
����]D��b�9q�2�*�_9����p�״�ǐo��f�� �>﹦WE])�כwi����CV��2���Zn��v�܁�̛�sqϭ����S��[kJ�۸�j�$e�/1p�+߽4K��g#�?�{�4n9����4~���d|��񊠸S�ߌ�����v[�Em�!q��٣r4���hJH�
����\�4�FA*�~����諢e{s?^*b�LW�zh�Eº*�^�'."5`܆.LO~ݙ]tL���LU���ĺ(WEO�1p�*b����Wn]��A����&W����L\)���M�WE[�b�PT���ٕ�WD��푴H����Nۄ1T
b�g���2<�}�{4n9��~ߦ�A�.?{3o~IK]*
$����w�Dʺi���Rv^_X/�W޷��2:ph�t�������dl��[E�\Cb�Xe��/�¾~ן�\*
����2�*�_9����1}�ۉtP�����i$�����F;�b�PT���2�~�E/�
��?^*b�LW��?	t\+����1p�*b�|����[Q�հmɕ�WU�W�~?�Cq�~���A�j�r"�x�� �X�P�����/�����T����2�*�^OL����q�\��x���1^��]
�|�L\*
����2�*�_9����1|���DԱ@pMɉtXWEO�ܘ�S1o��2�*�_{3o1p�+߽4K��];����XA�Z�j<k���{�v�śx6�Q�ƺ_Np\�k���EgRXՎ�1p�*b{���諢e|�b�.ů�nW�|.���옸S1}�_��5a���r]tL�����~T�Ҡ���~�WE_���
��'�n̮��T��2����ț��;���!���S����E�tT��ɋ�3��~��+�WD���~�T����[M�����"�fZ]
�|�L\*
���vetU�2�sM1T�� �Tt�%�E#�����4D�-(RPH,"ŦUU
��H�%�F�h��JB�����~��xXWE_h�-_�%ۑ۹hCrb�W���~�y����kա�n7�F��ퟄ�
�U�^~1p�*bo����V����@6:���ݷ&�9�c������Ƽ��9�;���E�]S������rW�i�*��LZ���]�S��&/Ԫ�n����s��WD��3�6ȭEq2��1p�+߽4K��]o�i��AS߷fWE]+�4�Ap�-�3Sp�ۍ�#rLK�º*~�����~�i��WD�ʅ�y�׊��S��g�.��tT���j�br�-;��� ���}�+�����i���S�������y'�B1A(3��f.�L[>7]��[���wۆWE]+ۙ����Sw�D�.�V�禍� �/�}���<��B*I�R<R���ˏU�$�I$� ����`-�����>���nx4nzO=S�x��f��ˌ\k��.�b�u�l.�������dkP6�[AY��b�l<!n]U*f��p�d��t�vƎ���b�cs�����`�X�lZ���䶝ʝ���9�pl.vӸ-�Aˈ�h��a�r!�G]���i������ں�c0'�c���t���e�뎋'ka'���[W]��B��p��ݳբlj闱�lk]��]��NX��ynjy�\k��V����߭�u���ؗEº*{��
b�-�7o+����홦*b�LZ���Z�q�a`fL�WE[�b�PT���ٕ�WDʷ���V�1^���t\+��^�4�H�b���
b�-��Օ�WD����3�UI#�A_�l�%�WE_���
��/��V�k�mGm6ܙ]tL�z{o`�S�۸�Eº*~�ɋ�1S����諢ej~2��)ƅr�1p�+�}4K��]�/�9��Ҡ�����2�*�V���*�p�/���$@El�um� �,��+g�㖁�P\�p���:i�n�3�	:;r�I 1ɉt\+��U����&.��L_�����!q��ޭCq�W}������=7���u%���C
��'��̮��C�K���H����n��(��@�d�u��t� �pXU�7���\)����K�º*~�ɋ�1S`��FƬ%�5r��諢ey���P\)���nR�WE[�b�PT���ٕ�WD�oK��#q+q��U���B��7q.�
��w&-���=߽�O ���}����9�῿~�ۻ���) m̥�p���ךb�PT����+�֫�B�鿯`�S翿b]�S�~N���f;p[�O
m���8�w�h��wmxw�Ԥ�C�8�ʷ$�rЮܜ])���{uetU�2��4�L\)���nR�WE_k�1p�*b�h�S]D��)#�I&WE]��ޭT��v:����A�dy����7�p���<���
Ĩ �4�
���m~nȭEqIn�p�L\�¿w�������a����h�rZ|��S�R8_Jk���4�e)Q��t�9�"ĸ�i7�70�����hX���,1�2�X�H$��)�C�1)7�(/"ڧh�hfF��bx��T\Bn�q��1C�TuQ�(dY���e �2��i)��,Ű�B��Kg����j���qȁ�vH�����:>)�p��g�g��M��<��f�7���D��	�x�PXY��JHQHD�����l�L��R��mM���/#[��� �-�5 �	 �
J�\�%@�2 ���]$(������bnlD�a��ki�����t�,Qt�Y�T�U�!�M�b�� �D�6��P:v��!� @������־�٧�y+�/m�.���M�Zw-�.^f������k4n7�埿{�M=��2��߯Ap�+�}�K��]?�z�����N��/
��'��2�*�^q{oAp�/}=��E
��w&.�LBپ	.�5.;��Ԣ[���.���u��e|�����`���Z��HZ�q��@���tU�1~Tl�߯At�+�����.�Wۓo
��'��2�*�^�^�j\Aˊ�jK�P\)��On%��U����rb�LTŻ���諢ey���P\)�W�h�k��6)����K��]}�6�p�*b{���ȟ�D$#R�
��G�V�!�L[鿱.��V�b�n�9-5-�G&.�L[�ެ���&W�ݼU+���NCq�+�7T��)~��(@ȸ�tj��������Ҡ�����M�AmF[��9&WE]+�/m�.ͤo�s�]?n����w�Օ�WDʿ����
��N�n;�N�u�)��Ά75����p��Om���gq�p���]��n*X��n�jb��۔�.�Wۓo
��'��]tL�8�����S���N�ء "�ĺ(WEO۹1p�*b���etU�2����.�o�)t\+����B����hdr�p�*b{�ٕ�WD���x��1{�ۉtP�����3�Ҡ�`���5a,�]�[�+������?��1_��]
��ɷ��AS��fWE])��F�q"@����.ž��K��tT��ɋ�\����i�B����49��Q�l �B��� �J�`Vu�
�
T��!A {�t�����~����  j��v�Z��Y��۽��@]F�=������n���U�����umLr���n����\�7a�s֣�;���΀��A2��cg��h�n+,�]����헿�~\��k�A&u;�9��'n��lR�z{Zv�t��ټ�:.�@��Y8���=�㎹ku�-�bڙv(xu8��fg�٧pq��Z��-��Y�y6���URT^@�+M[V�ݸ!2�1��Cv�F�zy}Ju�ݥ���Dڸ�O]�+"�����p�������p�*a��޽<��\~�>�h�P��r)T�-�~��|(WEO�-��m�r�U�f����=��O&�X��G���hr�¾���9ǐ{�g�F����
�5�K�"�8�%�tU�2���և!��;����C�I�9{Y�q�ȊP�?~��{����֮��u2�����p�P\=J��PO۳�]
��ɷ��ASۛ���WE�]lſ�Ap�/{L���ӹjX��1.�җ�D��ɋ�1S����+�������Ap�+�}4K��]?"��K�� I�s,Y�3׀��]z�&�\5���5���Xk�,�Ξm^����.�!rT}ߒ���߳���諢ey��U��n�}G�¾?f����f����w�WtaYxi�B���z�����ZtB��2�"0����H$�F�Z���������r~�]*
���?~����&W�7I� �.()/`�S�M�K��tT��ɋ�1S﷫+����󛷊��S�х�E�L�2`�Eº�~����~Ñ�߳��ӸF�;�`�C��{�(WEZ��i�\��-�$�������i�����ׯ߫C��n��?	t\+���&�.L]��a�Ah�k���v�y{�ɾ;<Y�G%�:�0ɝ�|v���ѧV����l<\&K~=�ʾ)鿮*�S�M�K��tT���
b�-�oVWE]+S^X�j�8ЮHܼU����.��tU���� ������諢e?ۊ�.����
w�v� "�ĺ(WEO۹1p���}�y
���y�V�!��+���.��tU�Պ���%��.C
�Sۛ���WD�~��U��n�]+���ܘ�S1z�j��X8ݻ����諢ey���P\)�/ۻ��.�W׹�.��.�{o+����_���mn<�.��u=���;�q�����ϵ�۵�y�^^^v�8j�v.�DGnܼU���ĺ&WEO۹1p�*b��oV&tU�B����.ſj�;�wq��R$�K��]}{�b��)��w�����!q�e{�hr��}��K�j��S��Z�+v˗ۓ
b�/���etU�2����.�{�M�WE_^昸V
����z�Q."X��;r^WE]��2���oAp�-��q.���S��L\)�����Օ�WD��L���Y�˷/`�U½�������$�4}��h�X*b��^WE])�_��T
b�^�{�/���HH�ۮf����9�c<�j×�����s�!���@L��zٹ��H��&ݹ�tL���n����ｽY]tL�ٻx��}�]
����հ���i����1p�1}�{o+��R�P�����.��w?b]+���5��PT���׶ܱ�ے۵.[�+����{7o`�S�4K��]}{�b�X*b����WE]+������Ȯ\�w%�.ž�n%�2�*ٳ^.L_}���諢e^���X.���=��8�b�ZfR�WD���M�������է�8�;�{+߫C��n��~�rA��"F>�ޝ��������?ye�?p U��d╪�(���q��yJ�;Y���D�����HsQ��C�)���d�B7Րǈ�c�4��U�{Rt��q��s����[���I���nW]�����W��}%ǆz&ţ��&��R�9is�1ւ��c[9.�r��sˎ^4t�b�T�U抆XԚn̙6�s���e�������-�k�a�]�v��+��hx��U�+��Y�s�rY3��۳��l����y(!3�IRv�.뻝zW���KM��r?����-����諢e_�=4:��p�{���D��#�?W��hܬ1y~_��ʶ��c��y]tL��~��P\)�}��K�etU�f�\*A�w��O!���d~,��rx��Y�GU��LW�zh�Eº*���b��~&C��է�y��+߫C��n�W�{ߤn��*���\�͇aq�U�~��.L_{�Օ�WDʿni��\I �w�D�.�W���3B�rڒ�l�\+L_}����WD�~��Cq�s��h9�!�P��_����T1uM���Ii�]�RӍ�\ʈ�c����/��+�\�n�Ŷy�ȼ�����q���+�W�e^���%���PW����]
�ԅ��b�X*b�����諢e7����E.۷/��n�{�N�F����7�q{}�Y]tL��昫����;�&J��`�Eº*���b�X*b��ݼ���&S��m�.����%�a]l��8��ˍ�.L^�sL���&V��1T
b��w)t\+���sL\+L[��z�Q."X��1��<��\o쯽Z��s��;��h9�V��,\*
����]tL�����豭n��Bf�4��gM��WEGGF���t�A9ݚ9טGoDI�mb�G+p�P\)���ܥ�p�����1p�?,L�{�����.7������p���i�Ev�;�s��������
��-���VWE]+^昪�1_ww)t_�]��U<j���ˈ�ț�.��/�o?]tL���*�����2)��B�\�B���E�tU�{ŋ�AS�=w�ܱ���v��"�諢ek��Ap�+���.��tU��i��`����i��WD����Gwd��.8b�.���w谮�~���V.�L[����&V��1T
b��[ۻ���FX��i�юR��v�qE����*��|�V��{\��gk��-�ahy�K��]}{�X�V
��Rw���i���~�_��n7�~���a]j��e�H��M��"�¸*b��z��*�Z�4�P\)����K��y��lѸ�QwC����.���N���WD�~�zb�.�����r� �{�4n;�p��{��A�.>Myba�b�%�b�.�}�ܣ��y��lѸ�Þ�~�y��.�Ҕ�ѠR�!#�
�<��x��P\)����ԇڒ��LK�º*7w�
ੋ����諡q��^���p�{��r� ���W�>���j=OI�����۬^��x� ���b��9�V��M��;v��[	Y�28b�°T���4�諢e?O=1T
b���ĺ,+��wx�p�
��x5^�b�#r]tL�{�b�.�}､�7A�{�4n:�p�ߦ�A�M��k�VD��vۆ*��L_?���E�tTn�.�S����諢ek��Ap�/}��ƙq���I���y��lѸ�Þ�~�y��ߧ����1|���]�V�n+	VX呢\�b�\1{}�2�*�Z�4�P\)���4K��]}{�X�V
�.����@�$ UP�v�Ł�D!����%	�@,)7͎�dE���`bf�.�ڰN��[�\��I�I10�j'&��4�	D$R_
��e�0E����i����j��r̓��$W ���m��dH��b����Q�b�qK�U�)ݹ/,@2L-�$���, �qԈF ����wI��@�             7m�m�     [@  ��        p  �l� h�!n�z�.Gkd�Y&֓�X�
�z�� �l���2v�F����Bmd^Xإ�K4���1�z��j�tao�Z DHN�k�mFE�ey�]�z^`+�Y��v��\��w*U��F�n�ݠⶫ�s���R$�iZL$��N��٧n�4����]s%�1�8�cm��W�dJkh�[s^VH$��a�e_UPnqw]�X&,$��2�UP彫��ػ�d��v��1[a�v`6.�6�
L�UhԫU*�Uմ]U�(%�3k�8 ����ol��ce�vW��l�⧵���E]PU�H�\յ��^6�v����H l�jiP
V����ۭ��U�'��X6
�ā����ѳ e���αA����V�۞�I$Zp9!��Ǫ�{n�cqT;d�j
ev��UX�	��mF�UQ�"�[,�
^(
�&�J����	�X
5N�kn��j�7�Kx)ԛKs��0�>Akv9�i�x��Q�N�j5M)��m&l9m虒�!dI���qOAQ��\(�b���⺞��6ztNK�M�%���$
�+����2��Vt]mT-��r=+��]���s�.a�U9�5��Dd��O/nɸmk��"�f�j45��\��e�Y;<�%��3=s��l��m��r<�nu���g�fKgʋ�]xr�x�!��a�c��'[��u�,�^kF"�z�W\�숲��.Q�ULxշ[ȼ���ց�u�lb��˺�
[]4�Gl!\�@R��Q4���Wj��]���:7al��ul�BC��v�ꦢ��m����ꄀ�vu�] q�l���5��b��(UUYF��T�-�\o��i&\R������zMoQwW!wyU���p
��WB ` �i��E"
�H�@�P�� ���6��U�(�D 4(��*��=����׿O���� �UԫU@U����=�:��MĽ؆�j��i��P�u�Gd�N<�NT���gqZݖ��%�AK[����3�7�H�'�ׄ��K�=;e�%��g�.������L^Ũ����3��F����G���e�ql��Ze&ufx�k� ;sri�Oh�C�}M�l<뭼�ݳgXA�Ͷz�$���x9z�x��h���>�G��]��zH��$Y����`���=da��͟G`�B�;�&�����U%�!��*�L�����P\)�����Eº*7w�
ੋ~�4�諢e}�1��rY"w��.�}ݚ%�p�����,\+L[���WE])�y銽I$�-t�/n�u9-7.!�L$�Cq��{f��pn�����<���n�*��LW�٢]
��yjl'."Ӗ67.�Z�
�syy]tL���*��LW�۸�Eº*7w�
੉馶=D�e�qڗv��WD��7oAp�bw�D�
�U����°T�߳�y]tL�����ܐ�e�2]�On��]�����v���9���۴�Y���1բ�ڐ58�o�z���a]｠�7A���h�w��ߦ�A�Z���.�����-pr �M^�A�n<����h���	�lGy��(

CjAn_>8T�~��Zy���s����7�w�����]j��e�H��Vո�ȱp�
����]tL�ٻx���?m��n<����h�u�ӧ�]�5�p����y]wԩZ�G<��P\)����!�����G��C���M<��\u5�,a��c��x���?m!����������>�����*�O��LU�޽��+*�%ԽU���u��3m���O��֞wg���9�8\&�ć,��\rb]
���,\+��/{��+����{7o`�S���.�W�S�Ū��5%��n,\+L_{=���WD�~�zb�.�}�w�WEF��b�\1z��{�we�rC+�����n�*��LW���Cp���$F� ٷs٣����i�ԏ:����E]��o�~"�$�M_�����s���7���n�u�IC� 6W�ZM�Y����$�lؕ��hRI*U���H!��q2$Ӗ��Itn5;�nn�=�Q۫v2;��X�"(�Υx@��h�^ �o=軺Q��Wi��m�F�_fG���7i�%��e���r6�������/Y��wt�wW�<�B�m�� f8�ޔl��dqo��wu.F�]� �&�&��P�M��|k�(^���$뗪"�����R�� ҁ�-V^D*
�EC�F����:�Ƈ��<N\-9ccqY���t��DD5��Bu���-�����$������w$���˖�a����a�\cl��i�������8�<cRw���:�VT²�.�����{�W?^�~�gU�k�-��6{]$��.��"I�Ce�"[1�>�wf�m�=�������>�<`�1�>��W�ّŽ�wR�z��^��Uγ<Cr)$�n9r.g�n�{�n柒���Fw}�J��aFC`J� �0�"Zl��\�SC�g��^���-�'����H/�W�7[#	$�I$�M hI&�N)Z��Vy���'^�����\�m�SOf��s�-�+��ֺ���
n��O<f���e9�lɵ��l��1��`٣^wm�Z���<�<����A�Q����y#7sc����Ц���Q.�m��gH�È��ă��rG�\�L�<�l�vk���3�xE��;/B������y�� ����t Z��㳼͡����n�^�&��rc��9Bm��W<V஧�y�l=�9	�S�B�e5|m�[��fhԹ�8�u�	�dL�M��P�̞��Zwu}D�Cﬣf�����acd$y[��wu.G���ߵ��w�l��}��	X� �d��{�PNf�
��ŋ��Vb��>G�A��2E
���z��۸�X��>������<�q���. �����7.��ό�lz�y�P��۱X�/�����gA�UC�I��� 
��ŋ��I 4V�Q�?o���wf���D��Ph�A��o[�{^�s�4�R�0#`r��`�;���\����~�o�ڬȢ�F� �g	��h6����6%�iZ۸�XO��Htk�P�D�SLI&���'u�hc�Ō;�$��Z�͍͓R�2	������}}��=ܢ�c|@6Y�bwu�V�G����>���<�vFgm���E��	��*��qv�<�oc���jNw��9[<�7:���@�o�H��ؗ����Xg��/�K��'��I��A!$e�?G�}3��!Zø�`f�)!�K�h�dT�R����6:>�����=�qz��<`�!E P�Q��d�V�k�(���<`�1�>�ޅhc�Ł�����Z����G��{�-��=2IH?44L_�#��Z�����w6j��2(�u���?�s��'#�{5��8x9�v�/!�R��$�\�[���9�-r5~?�����b^6��-���D#�}Չ:ļ`�Pm�Q��sf���"�}�^���1�7><n`O$��4�m	e��Xxڄ��	d�b��6�Z��\(�8�E��Ȣ_wW��r=ky����~�w��"]4JʊF1��B��������˴'e�.Eޮ����qB���WS�
��ŋo۶����K���4H��gc��$�9�'��;U�9�8�:�dm�1�����H�@՛�	e��XxځG�$���[�_$�8�C�� 4�6j��"ŀ�YI��՛��DF,<��L�(��j����޾���߅Չye5Z�Ȣ�F� �&I��x�m$mk���y�+BYn��6�$3|i!p����2�)6��_��٪�fE��}�g9�̿��W5���'������` ����x�*�Y6�����`{=D�M�+�P��,a�\�z݇��k�=�G����͍�NS�s�[K�pe��<��n��{nV���Om�v4͌snQ{fw!�ў���+f�!�&6�z�Ny�� ��|�l�\Q���l]����#��.n��:4H؞��K�#Z���;��Ӟ6�Y�G>�%�n�x�l	�68ݛ��9��~=�ww_G�}͒0�Evl����Y�[�EJe��oZ}ٳǫ`ޞ;��㛬��[�ω�-	g]_�<mE$��;�A�ܡZ���؂�L��O"�^���G�]_�K�iZ菾��]��^�2\�=� �a)��P�/�w6~����Z�ȢW�{���Me,�Cd�s+z�#�FHE"$(���{��Zǝ_�7�BI}<݅V2u3Q�����^��6j�ّįZ�u#����%洭�n��d�_ Q0����Lz�ݎه1�I+���C����j�A����@���;�(I-�]D/�w6j�ّ�s��Cq�bM���s�u�}�����0XV��AnH�X��蚎(�S� ��>�����Z�]_�7�BHlTnX��V"S/�6��_��l�M�#�>���O>�N�U�Ĩ�� ���3@���,�W���G�����!$4�xt ���P����@��b�ȣD�,įZ�u#ǩ��_���B�L�K���vۙ�1q׌���m�=����v8��vݫkm�7�O0�]��۱lK'mI�(�I-�]X���+A�wl���8孃�,y���E3=�uݚ�v���z�$���^Gu���(��1R���Z]�l���Do��#ԟ#�����WC�.���M��cTYFF��Ct�����$EּZ}�.���e�	{V�j�-���P�(�a��M��M(R�ڋ�J�!��PؘU�����T����[)旖h��a�.�ғ3_6sF���zt�\$�-&��34-\R��H+�Xd97�%&�W(�R�I�J�FHȱf�!�дiK�]i(�6�3���H���t�c c�m	���A6Q� �� P `�hl Рb!J���R�1@-qU���@<��V֑t��Z�z�kw9߽�o�ｕ$�𳉴D�g�����G�YF�T�28��a�@�dl��R@Vֺ�X��Ҵ%���a�j@o�sfˬ���0!�L�:�un۶���=i�1�s�ǭ��l^\s����`�L��c�TH�b^;r�a��QfƝ|@Vֺ��Ј�I����i��B�L�V�����V���(٩^"�@/b2 4(la�a$mk��G�G�#8�[5
�3�-)H\h�2��	O7u|ժ8�5Sl����3 �0��~�x���j��Me,�Bd��4��6%=iZ���XoZ���lt}�~����ܞx^��[���t]4�rܚ�GmxgU��h2�����8w��b�b��z���e��a�@`��͉OZV����$�$��_}����!$4��fĽ֡Z���aÍ`J� � 
�I!$ilwЌ�>̴%�꞊޻���vX��V BaĦ��^빳U6̎-}�n�_.TG�:��Td�H 	���	��_�tDGs�̿��~���{�Û��5�!;����n  6�V  u*�P���sy�ܘ�1�i�V.���s��#�����G��8�uͥq��G�܏]�nB���ǀ �ͺ����J��v\�N�icds�Ѷ��(	غ���\&����=����ݲ<�nW�{5ۜA����T�ێ��&[�7'$��C���)Y
�Zvͽ��{9�>�k;n��M�����jK�ʻUn��uշ�z8�gC��ɒ��Z�](�7�k���#��n�ps����,�[�BHٰ��]��Y���c)�A�h��Y%����V����V���,�}���"�.�H
��wPd�d� �c+5��'Ku~�X֡$>u�_}��$N��& 	=͚���͍�nR@`������3�7Ʀ@Q<,�m����޻���u�B�]͚��dqv;J�a����xL8�98��z�ݱƎ8ۍq�u��w=w_mg8Z�^& o �[-�7u/�*#���]�!:[���Z=ϔ$���OG�&	3PK@��Q�w7�3~t�28���wR�r�w��B"�x�A��,XCOwڇ;L�V�����V����lԯq �H�S ѡ@����}��C6l*{w}�s��D�p�!q�^��%<Ԇسb^�P�M�Y��Z���Q�ں��Z���NO޷l�j[1tG&���Չ4v#N����(^ղ��� l�T���'Ku~�޵	!�6,���p<S`��='��OٳU6̟�{NovBHtٱ��K�mN�ɩ�H�q?��fz+z�n���2?��w6j�ّ�r�T��i$IL�)����'׻��u�����T"�TU��߳~��s���"[���!{���ùB(f�(I�C�6
��$�mv�:��	ݰbCv����`(X�c4d5z���q�.z�M�OGfWe������M��q���w�^柼�P$��R��a7��Z]骁=(��&�4Y��Z��K�ʈ���w}�s��E�g�I��"�d����>��N�T�2��tDDDfa�b��1�T�ٱ���y	�~��۔�D@��> �dQ}�_$QK��� ����T����$���͛M���}�f��&����'�5����<��e��+��0��D�@m�&��H�321F�&�D�F{���C�"�}������28���T���,�2I0�6��?"#���ٞXd�p^���Բ"3�84�&�PhG���{]+Bs}>3T$��ś$T�3i"��B�{���OEo���_UfE��J�7��η�5~`�1����[�͌�j@d�śM�����_��@��$��WB����W����I$�@j� 5�m���7e�\v��A��s�6��9�`S�t���
�nkn�W:�vS�r�c'm�4�F�m�'Ci�r�ݘ�@%�X�%v�K��$�k�@
I��^�Vk�q�uS)vg�ͣsv������Gi�`l�vc�7A�b^�{7fg����b��Q/<Ri���m֜)��nq�c���ر����.����[���l>p�[Wh	��O^О��n��a���5箳'B2l(�y+.�D�26�(ˈr�.9}��������{]+Aֻ�^G[�	 Ȟ�4I3 ��f(Q5~���K�Hz���Dw[������aF�:��QL��+�I������͍�j@VSu~�����2�|� 6�7��Hm���S����#�s=������͎��#��B�EQS@��30��7�Z�^BC�/���K����l��+*+��+�1�+d���������x�n��.ݦ�Ğ'\s��l�8�lG�ҍ��=fG�[�����z!�/+�Z�p&���owڂ�����&"b����I�H:�9�bs�\��y�T	�F(@�4I�b͇��$�����ǭ�����z-c8�jLb �A��͛���ZZ�,��֡$�Ɗ��H��Ke�'�������_��e$o�ٱ�}G���L�@��p�{u���Ga�o$��A�)�q�O�ؓZ+�[��Wm��-����?^��csZ���9����V�כK�f�S (�4p6���mOD����T���!�t�f��Y�ſpʂ�x��M���9w]��o[����9�|,P+�Q�z)�(��a�"��S��o��n�}��9x�<���2Z-�C��5|z̎+�]��H�U�w��^0PMD,2AK�Hm���������6'3��Z���:ڻnv�[X�z�x
ۮ��ᮄ��� ��Nx�����^�v�.��u���Y��n����+xt߬ekiy	�=��*B�d�)��&�owU=�!�9��J���qf�f�	!�K�h�d���4��_�wڂ���g�o�W���i�.��#��lc8���{�ZZ�,��֡$ٹﾉ��}_v/!�/�&*	"	�`LUI_��e.��2_p^�;�}J�dklG��Ͱ&�nѸ�@v�9��/}�|vM�;�[rzJ����a�n�����˫\r�&�N0ɀc3 �æ͌�m/!!�/�\����	&g�}�ff�j�f�f�	 00��>��~�����]	�PP� ���H��~�7u���:��b~��N�\]�+��b8e�����$��Û62�����ؿX_o�jjbA��u�S=��u;5sV��}����9{:$C���J
�H,% Ă��A$E�����zY�eRH5JS#���dD1� ��E�T=�I��C��]�Z�	���>N�`���"QAV4Pޖ�E�|/r��h-KU�),e�H�Z;!#!z�G��v
Q
�*訑z�("��UB#VE'ÔR�J��#!�D$���N-BFA$����f��k�h�%�¯g8q�M���we�7�!�pڱH�)�``M��G ��
݀|Ď���8NE
�i�C �@@^��
���n��z`_g:�:c�P)Ԗ/х+9_>6�$��X�AjX���"���$B@����úh�����>���|��^BZ��gJ7E��'��m� ��             �`m�     [@  ���       8  �m��� P��������=t��:u�t��6Zp �m�e�F�qٱ�	=�/K��dd����V�t�YZ(��m�@<�t�<9������A/j���������:��FI�S8n֞we��.]�U[�:�v����2�V%�'�UCi����TqE�oP �T^�5Ӡ� 	���n�jL[@�t��ݶ�b� YTK:��z���.�ԧ2l[J�!u.��t�:y��/L�Q٭�����,�Wn�!6���a�ªڀ������
�U*�͢�����UJ�BXg����Z.�ֶxD��)�@j� 5ʵ:.�^YY�0�d���m�$��A"Sr4���m�Ac���� ݆�r���b�\���gN�Urj�B�r�U�z����<�QI� �R�����X :���6\jXȵl��Bk���S�VԺ)Y&S0� �Kx� 
h�[jv�k%�kze��-��̒��[Ӥ�a�a]��Qkq�r�u �=��ݤ�	8��^�!�l�-���r$�%���NX֜�6����§:��Ѷu�lӣVm3ԡ���uQ[/8�m��ݓu���.�ݫ�V�2�����m����a�g�KP9��눻nvywf��ml��'N̝� �jjbX��<M��֌��n���nsw��"�Rn��ʹ�ٞ�]�:�NY���p��i��{\�g�t�4�:+vPi)��o\���q̒�@�\;v�yw:[�a�Im��S��K��l��*�i�C�1
���ܦ2�� /.��ncg�zW���+\���;'UWv�$S�M��P�U��q��Kv�UlV5lJ���m�nٖ�kz0 �nW�E(�6�$jU*�S	����@�����Pl@��h��>M (,�t�ăa�[-"�n�{�{��w�Oλ�  �\��2�UU+��K��Лi�.�ۣt��+E�c�ܻ���U�B�Eܜ8z9���z�qk�uծGm�Ͱ@�#�6�Ġ:ov�73�ø�;��.6v�.^���N7\���n���0`vٹ�A��rt�v88��g���[��8۷+H��(��s;mtn�v�f݆헴���񑹊��ǡԅ����tj��vʶ;E�ьt����@V�sn�u�Q���yq�ok�ɰ����{�PV�//;q���xP���Ci��i�w}�+j��wu{��ϩ���4�hb+'`u��CHlY��5��sf�V��"#2>��U�{K |qA�j�K#�q���~}���g�}����Z��{�T�����m��K�U���w}�[fOE]�n����5��lK&g�}����Z��oZ�u/�TG�����\�Lz:�gu���v�Ü�ш��ի�z�1��h8�iz��lu]l;K�4ߟϐ�����?7I!8u��ĭ�t�/��-6����K���������UJUkt��t�J-ڡ+^|q�������{�f�2z%��T���xS-�H�����g�޴��κ��oZ�usC)�����jh� �6o��s��Bw���c7Ν�B��z+��I/cķ͇�{�ZYbŎ��>���s0:lؖ��}}���l�a�BșnB
�%�gOc�x}�u�^瓪A7;e�cl���[���qͥ��ha)���]}����3�w��o��Θ�ܹ�-(��hSL�����ݚ��̞����wWa���8;Cr_?UUUW;���}�_�d�[� ���$EB�����/���o��bv%�	�2P��IJ�}k{�/X�ς]��wR����[��hm��tH� TI0h�,����s08tٴ:�ݚ��̞�oP+`2�	g�8��8!�G'{\��p�]������24t//�oOL~X�0�;��_Q=��V�0����Y������b��1�Pm1C�]٨}l��Z�uq��8�i����ЃH��ZCb́���ԹUDqSz��W�P Q<h�p�DH$����Ci�͛��
�}��|0ś�0ģ$�5UD�$R]}�,��Fľ|��ņw���cN������h�xn������m�n[lIܐ��v��gBL��vh�5*�ޅ�9�պ8J���(�,��#X�`f6"#3��b͎s";��$	C� �hN7q~����$6��ٱ8^��������Pȫ�0jA i�qI ��;�!��`B{���`)ن���D�DI��Y�8�������Ł��I*��m�0Al�Ȣ���Z���s8��{o���ٯ����B��%BQT�`�@##P%%#	�Y��GO�o�  u*�P���]d5s���aF��{M׶(�6A��ݵA�N{����ǳ`�a�Ŭ�/%�^{p�w@o��:��"\����;m�(�㮽v����J8��d��9��r����Y(N����Z�sűV�l��dճ��U�@��^�mF�M���:��d��Dq��θ�p��wi���ۮ����PNy���ߟ{��o��%��qy��,�[ر�6����U[!;�N��}�pWk���\����|L����ߏU���/{�,��_L_�DD"�s<�C�_\�H�`1T	1~���t�菣0�q�b�����Cw�Ջ���e
�DMM�Nfc�1b��wujٓ�}��wuv��$02` /�#�����.�h7��b�׬���U*��g?����~w�&�A˶�)%�q~���u��٘Y�͉�wҭY�*�߿UV���2̺*��=���`z����*�n�`���e9���6��;
n��"�I��4��7��z<�,X{����bH��k�M~��z�����-~n	�!r;��z��璥���,T�iJ�7|]X�1�(�$M|��X��#��Ȣ����
�3�}�nR\_�pF�o4Lɐ	�`A3D��V�=e$�9��i@
'��'A��_wJ7usV��^�l���LQ+�@x���8V'��ݺ���v��g�;��b۳�h�E�z�\��ƈ��s���o o$���u^^�"��;��
�3�}�(���`��M`x�2hE�}���y�k�%!��=e$�/Q�Eh*�@4��Z��z���~�~�埏�աM�.U���H�ZRv�Yj��D��m�
���w���n����.���@�>C�!�i��_^�wU��2���l�`^�]��^�2\��Q�61"[���Tq�]͚���%���uv~�D�#l0��)��4�x:;p0��vܕ�S��e�v��hgp`���][�[ �L[ēW��ըWi����F�j�W>��x��[�ǒ��Z�.� �^�wa��Ў�itx��n<8�,lbl�E��7usV����9u�٫�z��ܹA�,���A��u^^�"����B�L���J˪�T��s�;��k�xȁ�K���"͉ǭB�7G�ذ1�RA��o�[{wxH���2�j6AIm�d�<�fݺ�y��gGS��]�����v�/�r�Y��H% ���_�f�I!�g�����}���ӟ|:$���Q&d�H3b���]�Fa�/�,X�g�K-�����6����X2�Hw�~�u�q�o���)*���]��K�k�ԏ�h�1<�q ���N�B�L�_wJ7u.V��WYlo ��6j�^�(��vw�{�.>=��{���qR�UU��P?t�z�O'wi������  n��^���6Y׫��8��0��=��`Sn ��p9�V����kZ��v�gx}s����,�\[�������7�[�=�����ݻj,���y���y��۴}��̰��E�Fg�:�ە�Iz�x��ZbĬ�6rI=�P�u�hp���,@�K��b�M�.Pp�FǲYfj���r;�nM��d�ֻ]e+<\�,�=��{Ƥq:nM�vv�s�q�3ɼQ��u��x_@<�ݫXt;�t��k͊3 �j��P�A�����I 06w������A{�ڨ{ٿӗ���C��<�l�S,2���yz��+�;��ޢz/��S����sؚ`��E7f��֡Z��lWD�;��Ǻbō�k�0�]����_R��_s��RH�6'^�
���+�~d �E�_[w7u^^�"��;��
�������m��C a�� 2
�7i6�cl��v�-���v���q�9�ϣ�Η\Ҳ��m��~��D:��٫�z��_[w7uV�h�)�x�c"��KIG�}κ�X���IXٿX˝q>a�K|��^�l��v���۹�߾|�������T��L4p(� W�ȏ�;�]$��l߬Kz�+K��1Ź�ԭ`D�0�4�n����͋t��κ�X�����3�}�����?��;;��ᝆ�6иz�ѹ;�-��vD@����\
���u�,q�
%y	��ZE��c5�~��k��'��@�I�j�I ��κ�X���IF�fķ�B�2����I�� E#��8���W{���-8��R
^��D!QOX�M���]=�c��C]�]���-5 򑈚0��7l��, � �}N�� b��ض�(�j���ő	 �R@`;)`�
eDi�$J¬2$�in!�ܑԉ$Ch�!&V!Q�$E2�&������	R��8b��0�"�a �n�8ܬZ�i����X�ceD ���>��A\ l��M�-Gmz:��J�z��"��B �m� Y�""�Q����7���>�z��������33S"L�$�ItA����B�_���e��ύc'��������T���E�{���Z꣊�v�H!�����&��n�-�.ǭמ��Ϯn{uF�'lth�g3��1#GV�[�f`����_�#��]��DQ^�wV�U ������fz.��N�ϻ�=�6'��he7qf�c�bQ�4`���h� ��>�-���;Y���z/��S�����	�F7���Efķ�B�2���c5۔���1��}P�$�w��q�����L�-@N� ���X��"7m�f`�5�6%���5^��$�L�� �2�`��B$�t6�'r��p;v�;�u��n��w;tr1s�]�C�!�I�q}�Q�����W�wO���F���g�Z($vV�L���
M��F�fķ�B�2���c5۔��&$�<0Am%���s��P��3�^�F��U[�n#���l3�o���B�2���c5۔��0�Y���k�g�W��&�E�	&g��ҍ�U��8�u��5|m�]�{��[m�����6ݛl�q�GN*�ݔ܂恎�O=s�)w`oS�q����E��4K]���usuۣ�Lk&��k���bȉľ�(]*7l�挴�N}%�Pm:��:i�'"N�d�|h�vy��V��p�w��j87X��۫����.�/]����F�:���Ny�g���7Ƨ�Ӱ�Y35f���p�#�֍��C/i�g��p��0��w;U_*B�$�fr��I����q^d�\G:W��uŌp혶�s�9*�nQ'Z�]x�g��t����v�wU��Z^Bp����nRC"�v�x�8�"�Q�;��٫�l�����wW��{=�ƥsx�L����/!:[����nR����=��#bu�(W��G����,`���G��7u|^Zc�����P��3�o�@₯  �@6��_S[���߰�R���6̏�w�ӽ�~ݶ�!�ԸZ�@�j �l���{/iq�S��lsx8��,��1��C�D��/�.?[��C�S=�n�uQ�םgO��	%��׽�hP�C���"�A:"�H���k~��/���M����w��UK�I.���X�.]��n�XM�JH25�&">��js�w��;�#a���(Ě0MT�4A�e$2���8���wڇ>�z+�J7uw sՀZxB��H"��.?YF�W�ّ�{���=�8���'	����0��8 �U��8�[qlm�p��ۭ�ټ�����m�)�0 ���owڇ>�z+�J7uV������o�/��ĀD�1� ��⻶�d}?}��:l���(N�w�ԕW;U)�����n[�-7!�{��������ߧ5�r+"8(P�J���>�ޮ�=��ӽ��7 ���nD�3SD�B�b;���]_�k�r�U|�-�Þx��G|�i�o�|m�W�Q�����#���u�W�?ͫ��y�f�[�#m��怷c�a����prЫ60��Ny�u�6����V?Eץ���TQq��7ھ6̎.ϳ�}�wrY$;���UJ���~;8��|�Bt����A�k�1��q� �"�d�H�D�b��;r��Swz!mt����/�'�o�7NBF��;��J ��]/Xom�H25�70B�}��Xh���3�0Ri�� �%��l XhK%H��(K �KWv�KZ�ha�)Q�*���O߯�׷�?+�B�R)-��+�(����e��u�z�>�z%۶�d�[�5�e����{Ʌ�������:;lY�v;Pn�`��^�����p�m��U��8���N�W�ّ�{����9�%�����Ȣ����P箯�7]�It�}�E�<j	��� �"�����a��$�h�acwuj�i�Z���M�軬�R�bō��t��>���:;�#c_uD�h^0�)�Sy���^�"�~��C��|�?{y�{���]^�EP��J�ڰ-��A�D�(���а�b�LH�(�ZR�E�b�
�T��� 4�B�c&#
��,Z��cƆ��(F5L�F-2� ���,�T
�!��l"	�TD��X،YA�H�E3 "@V0�R4����z�������� 	�m���ո�%�h��1������Dx������|}�y��յ1�dݝ�*��p=�B�r! �w.9�[@o����\-����+-�4Nl��S�������6�L��!�眇+�8S��xz�1��u^3":��tң	t�y/��Y���]�1bH�L�P�u8�C�v-����iko=I�yWqӰQ�/VRI	$[�N�:�<F7
c�֛�{n��;t��� yO]�[��b��w��Qd�.9M\��ۏ����}ο��#��w37u}��dQ}�9b �&��Z�>�z.�(��_:���޴�/��X��ǈcH$�8��swWܽFE�]�Z�>�z%i �ҋ(,a��67uWΨ����;�_fG��n��h�� �c"�c- ���W��n�A�,X�Q��3�o�����ں�I�3��m�txB'Es&������H��k���9O�S��8�ܜu:A�h��&ߎ�W�ّ�m������2�����0 �_\� �	�bO�D�X��{�Ο{�7��.�XQI($c*Q�0jSt�Q��60`}��s������ޮk��l�����Zŀ�%6Io7u}��bŅ�����o��}Չ:�D̘�(�,X��vDG��r�6;��w��Dfa�=�,N��q�L��������z.�ZwuW]QE�/[}�n�ka�An@ Ԁ�㖯g�C��ɒ��cu��..n�Q�#I��.F�Z�\�Tf&	 �,6ڄ��s,,e�
}�dǵ46��(X2��}�(�]_A��_u"��w,6ڄ�Q���.bD6Kc"�~��C�����T
�.$�BS����z�zk����y�V0ch���Ưyi��Y�V۹���z��-����q��DD��p��<%��X��!���Dw_��A�pE�xr��RJm߃S��b���#r�mۗx�.��v�!����u��וxƹ6pJvk�la�S$��wWr�[�wuj}D�]޴����=P%���e�
L�}�XE�~�����GwvFfǺbŌɑi��0V�7$���=��3�����R��x>�gOqE��LЁ���]��M���FH� �1Q��5��~�������w��}��/�XR��U$=�9�ov�/S��r��P	4��b͍����7]�n�6ڄ�/��6��6��<�"[��$��l����d�3�VS;	�[�j%���p��`��)��-�u�z�_Q=}�N��U[�n#�<�h3��	����g�1[n���g�ߗ]׫��P��A�X�Sbz.�֝�U��8���H�k���>�V��`-	M�����3f�a��E��}}+�=�u$��H��� <!`%�=�i�j��	|{7��޿y拏�V��}��N�[�Hjm�f�@�~�;���"Hʔ;�3�H��O�hNC|����-#��VP��"�Il�
-`WB0ʙXCBD�CF��s�<7�С��/�4r$���)�r�`�)� ��o�^ek��K��L'hx��)6Z���4�	�j�L��N��G2���"#Qx���&I*�d:�C(�l�"d�A�3�%.��(3�w�w�d�����X�ې����Ӄ�Nҥ�s��QEnH�p�G��C�1�X��e��tgFD�b��W������h��$����s3333������           ����`     m�  m� �>      �$  ��ۜ 	�5�ؼ����g��wb۲6����]6p �d�t���ˬ��G$�)!i5��V�e�S�n���g�-�m��_��˺i4��P�h,�[P[J�T�J���n��hj��U/N���rv]��ݰ�����L� ����7Sq��*�mm:1�ݺ��=���U��&8����^]�N�r�yf6*GJ��d��#T�����3ڍLK\�*�U"p����ËhW�Xl5�G �pU�)-UUm��v�^/ e�
�݇j�d
�
��!pr���S\$kj3���t�5Y��H\յF��U�j���g��������P/l	i䒥.:^��E� +�ŕ��0۳v_=�0P]<q=�2ۉ�:��b��=Ml��+U�m���U�[S�(�Wnkj���V�Mm�n��m��ѐ��
7j�
��,��t�nQ��p$�N��#j�A�����$�6�d���1�[j� ��)�to���})&�.��!q�<�����3\�`BZ�s��Y����Eت���]�M5m�U�8ẞ�7J/h�):⪐��n��,�R�Ά�זtf褅]S�\�ZyN���}��.ՎӞu6��&���v����=j�v��5K�9��H%�tz۠�6Ӧ�3$�bI0�Wd�ۧ�#��k`�{ܫ�8���xb]�^yM	�tW\�Z�"yh����C0�%��M�T����xӔ1Ń+UV;gF�x^@X{c#e��5[+ذ�1�V��t0Y�D���2�K-���fc�C�s�(�X5FĕԵ��;��ojUT��b�p�8(��F�Tݴ��n�4�[WJ��DH��}u�M�l�M� �[�-��q$ҵ�v� ��/A� ��Z�dn���UJ��P�U���S��a�(�[�R ��!� �&P V� S�)�+W*Vw33333333�}���J�qJ�T�,n8��@�պ�Nغ�K�hSn�F$�$�HsuN��]�G]�']�e�����r�;�T.�ɇn3���i톺�۲ZM]�]������%��`	��d*-1n�ۣY봕�Z@����U��K����&���
�f�iҌ�.�C,i�p��glv�u�S�!u�����nnpE�6���E���R�`��*��E(�Iݳ�q�;�Ǝ��r���bm])pRr�-k���З=v���Z��k�������M��盤����}�[��^C�ϠO���m���*�U���z��/�]w^���OEq�<�U�,@&�H
�f�bw<�+ﾈ�=ܽ*�q��$�ώqŉ~B�Ka��q}����������wR?us�w�9+1�H��Q�}J�mߥ �.�I��E��_$�}�G�z�%�c��L���B��x����l��=�m�����5s����ɦ$�MQ�"j���u�JH
�f�bq��SU�xC�i���-<`��kwR��ޭ�N�Yd�RB����xkH�8���c7m���î&�MQ�h�B�&�bw��J�mߦ�>��"~�-�K�����D ���Ïi=E	��7��nR@Vk7���Ҵ�xX��ǈcH��1Wz��K�*#��]רu��}���� X�@➽�w�뱞�Ve���^z��6�M�9n�J˫u�H YE��67u/��_����u�n�q��$0��L�@�4LUP4 3f�`֒��H�}}+�kwҒK�u�� y�h$�~O����U������=�������0^e}_�qw.��Wޡ�ă(�?����Y�nR@f�lX�nܫY�DAl��63�Zŀ�%6Jl����=��3�i}�pK/��c7m�HtE>�&x�?I�޸��4�vv���9xN��K�%p���竊�.(�q8�X�G'x����]*��qb�8�I	Ӳ��aE=f �&A��3$�Bt����Ik�Q|z�7��d���J		�%���a�l$���s~؏���k���S=ǔ�(׌�qS��u�n�'3����;�_���g����pBT�@$$DAdX��"�ITy�ߟ{��m�Zj�����.@�Ս��"�}�G�����}ܡ$���?�����ڎ}:�^�qld8ojwoX��� ��s�%ի��y�vyzM�v��ƈ�T/ �w,3����s,nk^�6�D��Ɩ^4
l�E����K�������j�Y�E�Zp-x�Od��5���z��.�u�z�>�z.��n����H%����)�1��͚��fEZ�uw/Q�E��D ���A�"�G�G�S��^A�r��^�u���Û�,aN�?(- T�$B�YZ$H®��,`6@��ەW�%,�H0K�����^���� j������[U�Ż ��܁�@�NAݰ�6�Kv��]��{�Q�5ӏ9Q���x ��k%�"um�n��x}��3���햤��p�klv�!��4g���ݼ8�8�팚wv-V�<����/\\��>���Dv6ZӬv2��B[�ɸ��;[���g�qp� ��qŵu礶1��q��2v�s�rU�fed�&J� (T���$:D��6l��9�u�nG]�r�q�.�s�*Wi�J���C�:�d�a琻�w*��?>����<�?fO�1f��ֻ�RK�8l�����~���22\C���f@=~7]��}�ovFyc�,Xg
����C<kE��V<%[]��Н:��Ⱦ��Ā��7V3!�S�0	 �:���߳}��VdQW��wW�
�O�Oo{:�g�H�4��4J.9|��P��񺰩�P��hw,w����e�,cCW���,hf�g��u�x����]����wV�^e�ɘ�$��]���6?>���ݙ���Xw������� <!`M7Zm�9H	�	D�6Oܯ�U�j��ǽ�G�KbhaG`6����ϩ��޻�����Zm���_IB�K,�,`ĊO"�����\{�Dq��٨s�g��yO"�x���3�&�n�W��1i��o�}�̊*��u#h�1��%�xq4�8��dsp���/��&�Ƿ`�k��^U3������y��/�-����}L�V���Ծ����$V00�#e����a�X��k	!���6lf2�k&&F��[fz.�w7u/�����@�@"4#�"��j�"�(](: b�D�dϽ���"��Ӂk�Zx�$�q�%%���J67GrE	Ӯ��ǵ�FbďuL� �4(H$�XL6�1�qb�Y�����ٱ�}��L��v��1�j͝�8f����ш��7d���s;�������v��c7�>q-~�W�_U���j@c~'��U6�/ 6���=��i�Eߺ��\{�Dq|~�wڇ>�z.|8�T��x0�}4$���n�*m�^Cw,���|��kE��V<%^1C~�v�ܞ׿W5�W���~��s��I�PA�@QqH�9^����w�Ox��!�l0�~^~�����"�oֽ�C疙��n��ܼ��(���x�ѝ�Y�����n���'U��;��q�u��Q��1P $D���5~��Z��ߏ}��}#�����qb�Fk�
d�0$T�A���0�_�J�Ҵ%���a��WR�K崙��~N�h��������c��D}���	��~����XC
82���+��E~빻�}o�1i��o�|X� ���P,X)tDDD}�w��K�'7�+B}��o[��ޔ��UAEU4�	/�'N�������ߠ � T�J�UҬ���{�_���6��i`�w6�.8�<g֕����gI�v��nަ:�i��@"��Zݬl]���M�1�'��6h���V^�K�戲���;s��sg��,�M�u�ds�Sn[�����Y�3�*��n��.I�������˳�J�ɵ�96�\���'��4�A�;g�Z����y��i������({ԛ̓2��U��ޗQ�#�;u���^�x���ޒ���e����W:p�DP�~5Rd�@� ����7V6�o�}�̊%�Z�u0gv#�.aD�� ��Ĭm+��BYn��kP�����Ċ��F&�I=����Y�D��{���������]UdA�-~	�h&ٞ���n�W��1|o]����Y�E�i^"��-2ZI��\^Zc�o[�5�S=�(������	���_�n��>��nZ
�u�Rtݖ:��t�t�ԇ����ڍ٣`�稄r���?����f¬ۋ6�g�"G(�uf�9�S5?��mTƦ^g9�\�}��&�*(b�I$W�� Dl"!(�WA ȋ)pE��ɵP ,�-n�H�͋�Z�ńk���$Tz �� H-}�s��I��fĭm)�|�����Ra�X��M��Kfŉ�mB�2��Y���)!�L:d[.A�]��%�q��UW�o����~��^A뾔�������ꨓ&hQ"�R$n���+WK�i����Ǻ�Wg��eG�.
�_��Z!���	[�/y�6j���_}n���W�w�xqbaV����m�IXٿX���/!����]�u´����a��wW�Lqw�s��NU�ѮP���)F��+�j4h[�B� iH�����p`lS�|͸��H$���
��]X�CrФ�FB�Ɂ �A5J3P	!��@�d�B�T4�R��$�PC~@����[�������mc��q-#�[I�Qb��5CVF}c��E��5h��w�*Ē�ٙ�8c��Բ�0̢�!�J7�HHH@nHC(i�:+F�a�r1���p�n�#݈�1]�6D� Q+d�"��Wj^P���T�����+�.s���6��v�=Qp 
 �A04��"9n�����B �I�su�~Py���N$6*eǺA�dLɊ��"͍�֡y��,��mBHa�Y��\������Ovj>�z-��7u#��g?UM~��/�������]F�j\�/kn;tl��wOrD�=�X��9�8��mt��#�@0Z�1$S��_}k���B�B��vj>�z-�I�Q��$0���ln�+7�Y�B�Z�,�����11��%��Q-�1�/�wf���g�߬�wR?Z��$\`6��(���s����D��	J�%D�k߶4�ϊHa�Y���}��M<�j����"�k�L��M�=�e����~��Dk/�0��:�ņr�̘&bM�y��ݺN�d�qL���ݟ1��DX��b�q�؈��0�!7���Kl�M���慦;���	î�����JHnďK��'�e�JI����]�z�+2(��׻���m���:��İ�P��;�ar}�>��_�-mBH
����ѭB(�p*��"�� U,X)!Ѿ2��Bs{��'��XӕLE9�L��L�P �H
����ѭB(n�qb�x�I�`�$��]
˕����W�  m�`m�^��
V���˺�����c;�"Nˋ�vΎ��n�z�pk�;�NӋ��b��d��H��[H����y��s����[�ݩt�uA��g��s=���ݗ�����O��ݓr��6[Z)˞��m�aw]��[n�NE��v��8yb��[��mӥv(��Y��항t�]�#���m�Ж�q���vn�ԯn�����wv�{���O�M�U\����yz^p0���Cjy���4on��v�؀�@j��F�a����5�_>JМ:��akj@Sm�E�~���`[�/y�5�Y�X)!�N��bV6��ώ�w�b�&�?H ���}�A�سah֡�VdQ}�[�h	a/�d���ufĬm+Bp�����I����HL0!b)5[ˮ�V�2(��ҒD���㎮��I1S�D��������]�6�ד�6{��h�mv��G#��Mg��bhaG`$[�f������z���V=��RT�s��{����n������]�����{8�$�b���"�QZ4��DA���D�p��.��1��A "#���/�͉��JМ�9�XPr�f�0j(њ�d	 �lY��kP����?g�v���%oW��!�>��Ds%�RMY�}���hN��akjC_�1E���/牡���I=�z����[a$
�VlJ�iZ�~��H9�����r�<���^mΌ'@K�c�`q���gU�gP/a���1��������?������[W]�z��fE�$�q	�  ԙ$��)��Fs]�hNL�]��������%���!�1K��p�r���f�E!�Tm����j�Թ�8��G_�
��JV��5����}��Ӊ�=V,c�kԾ�2Z����"�O!�m���\��8���vj;L�W�7I8�,��g�������l&;l��\]�c#����x��$�Zi�Z�B!�B�Wr�_��1��"�6n.��)!�K�RE&��S��f8���vj;L�]lӽ����窕T�zůQq�." ��G�Њ��X�l���e�%f��?��-�R1Kh�(rK�s�U%7���>�����ջ����p�s���H`�eB�
1���@��$�DR@p�����wf���E����W��I�W�gy�\R��vkиz����A`�W*��r�\	��[\ٌ�Fz�?�a���ŋ=g�#3���Ň_�0&�pE�٨|�3�u�swW_:b���j��c� P�B@1b�OYI��,J�iZ���Z���Y!�H�&�n��Ϭ�:�Z�P���X�l������"�T8���L1C���B�L�]������=[�؜��@�� ��'��w��������  5V ��Z�y�6�{���*��5�[t����%���rk�GS�5ӏ9S��[�vp7��nJr�m�VY����wͺ��09��7��b��������>�h۷9@@��tg���|�x�!�g�n]�c���p)�R8�[�'�㭗�i[���t_,��q��=�6��l�ݢ7�=�������n�g���g��7��U]���Y3-�� |8�nZ�).ǭ�>�{z��TmRv�]=l��8�=c�$�A�_ ML�}�:�ŀ�e$6��#�}�]٪�V�%$0��l&���w�ICbͅ��!�;�ڪ��E�)�F&�����8��uݚ�v���w7u}���K��x�$���>�����|:�ŀ�e%���u�?����؏����.�nw��67W���IF�f��Z�mѸ��N��Ef����L�k��x�yɸ۷Y}���ջ��w;u�#tG-���V���VޯwW�C~�5
�3�s�\8t�C�-4ۋ���������@U����}�D��@�-Ga��uŋ9�I~�������܅� A�7��}����,�W���IF�f�11�IYx����٫WUfE�����ޣ#�o�wf�G{ō�����fz.��$�D}�/�(f��!�;�7t�\o��q]�q����.y�X���=yC
�u���Z���4WjL��	)!�\��bVkJЖu�DE���j��;=BxSg D,I6c�~��j���d1-�^�.�'��}������H��5
����w7r�a?��0!P��(R E��id" 0T@��g�[��;��_/���s�J@0Z�1 S�b[z��\]Gߺ����~���g�<Y�������rC���f��Z����Հ���[��vڻ;g��u�3�pu�l�w.i1�I�j��{^�x��tfu�p<!v`Gߺ��B��z.����T�Q{�����.��K�W__۳���*����$��6%f��>�Xy� )���Q�"h�W�{�$���=|��}���7V1�SP��L��L�P$��Dr���V���_���DG�T��*��w����ᨻ���;��ٛ62���cf���Y����r�͌�� ���u��==�]� �U�n�(�m��9��no)�y�a��7e����JЖ[�����$���62��}xF�
ꊑFf(�Q�]X��qtQC~�5
�3�s�\8h	��&8�$�wU=�#������_Z�C���usW!���ĀE�#�,֕�,�W���I���o�ٱ�Lk�Ah��<_��߳}��\�b�޵��n_���W9���o��?��m��P 
��  ���O��ւ*?땭k!������_����QQPJ���p������DDDD����O�����?�_�_�����^���g���c�����O����������������� ����������� �P !�������������3�p�� ����;������������y���(�����Q�� �D�D�DRE@RQ!H�H#H+H"��1D��DR
�D�H�IED�Q ,"�H��Q"��D�, T�E)H�E*�H��AD�D�H	H�H0��RH�D�1D��@R(�D�D�@P�@R�D�!H@R$Q 0�H*�D�H�$Q""��	H � �Q"�D�H
�Q"H+HD�HQ"EEE @R)H(���E(�E*�H"�H�� �1D��  E �H"�"�AC��(��H��"Q" 1D�
 E �EDR	H�Q 	HH!H�1D�
�Q""H 0D�	H $ �Q"H	HH��*E(���D��"�H��E(�1T���E������� C������'?ȳ��� ��m�����G�3��/��� �W��!����a����ߨ@ ?��� ���?��~� �:Z � t�/��į�0�u\?�U��?9��j` � O�������?��( ��������?���R�� W��j�� q����H����EW������9����  ����{�H���������  ����W%k��B S������e�����
�2���|{��� ���y�?������ @�UU)@��Xh   (   � ` �   z            dUU U  <( PA��f�UG�m��z��d
;���Gu��f
ic��l=�̎CM���t��ݝ�z��@����P4trӂ��F�;���|�"��N���ԫ�m��rh�rzj��OC���S�fG {0�=�O��	�����>�h�$|���	�ʅ _x�U<tdN����<87UUk�w�n�P2�U7tjΠݎ��j�^��I�US:����j�����UUv�&t���T{{�6��z��UK0eР��Y��_Clyd/p�vUs1U�ݕ���E��	ހ���ӻnùҗn�CM���h��t:4��x�C���kxK�ѧv:t0���`�����x(�ɧCN�����z2r5���}�����龄���:t(X+�c��>�E�@��+A� 
   � �D�*mL��!�CM00�~=U*���j` 0 �ɦ�� ��U*FU2 �     j~�T�P 4     
H�51'�zI��F4��F�0��!IU!�      ;�����OO_�m���DCN��DCJ
���(�y���*�O��J�F1AEB4%-�REDT��QBP�HY��F4FeP�Q@�He�NH� ffFAXe��4%�DI�e���E4��Q�8A�e��AY+�4a#CH��Y�T	��"!��' ���1����B'�ED' �?��{���Bk0(Q�  ���������>?,r�sW��F��f�+sc��#?��Z�ڣd
:B�L�2r#�f�h�=�SM�	
��iRRKQQ�ų0��]6y��]uN��r��ٍ�3Z}������ҕvSΫؘ�U��bMYA�Xվ;(R����˸�����j��¶�jC����[���׿v*�EC$hW%�]H�x�@�D���P� $ 7= = �
Q�Aw��
;ș#�(n �AC�P�@7@CR��@9��	�
s
�j@. ��qGP��@�P9�҉B�y��C� �.( D_DC�(nA�@Ԡo �0��q �@��!�P7��"���AC"���\=Ȇ�!J�B���;@�� j8��!�q ��!Q � 7 �C"!� d d�o�#@��C��q(B�!��m�	Ġd�R��@�5(BH���
28��%��
)@ԡ�Ġw�@�0!� w���@�ԧ� �Tu��@u7�Ƞv@Ƞ\P;�B�aC��D:�:�9�N�C%� �P;@P��9�����ࣨ"� �h � H��:�
P6�� � v�%��C�y�+� v�
�;ʹ�s�!� d v�J(�� w�
U�I��P��D( ��0!��v���DW �H"��B!J�o(�@���{��9�[��x��S�,�����\_�K�?�"~"�?��'�W��R����'ܐ�M���+bfX�vk���X�6�&D�)������wb��e��me����s���!�R�	�8��4��Uͮ
�u.nNg0ff����A#��@�|A�u"��d�$x2�T$dy&�Y�d�]tL�yJ��4ֳE�Ub�f��b��.���#BӅ	�X�U��1z�C�uU�YT����H�`b_hN�
E���6޳J�C�BEtlCD˂郱T�i�5��#IG$�ewYy^�3�������>�an�m"0���bq�%�$2H���^����s�Mʭ9d��!��1�.Wk�"m6H$h�Vp�t���ۂ7�E#� \"4�`ї3��,%<����+�H=`xLẁ��7�AlC�A��mo��ƅ��s���4@�@��:����r�kvm6��e�=]*L�@"�×]޹/G�C��5&�B�ДY����] BG�x�h�P�:�wǴh�u-0�W�W���s��+�Cy���=���Sޔ�S�zgM%���p:Id/��«!����b����BD��z��G��}���3�ruz� �a�"8ú..t���L�,��:�!]6�F5���
��8i��ŋ��H�
B�D��>�V�~M�� ��@v��SJA���' ���=b��z;�H�M��6�a��4�=�ӷfV�xZ
�V�,"���P14`D*!��z:=3|!O|��c�C���p�tm��	 1H�Ƌ��a�I��0�F�=8�
@<��h4'+�%-�6�B@4hm�mv�q�`Xʹ�,=�aA��ѳ���
[����\�1�3`��'�&�3�R��{�b��@�9�"��,*ģe��Db��]h�bۣn�@��c�n5�vq��M�B"�6�8_n�G��A�B���#���T�^��<)��JF&�D<�@�,�Mt�C���R�a��HN��*{��w��X����5�)��A�fw���#��#��^�!J�;/�� ���h��B�䮇B�%v_/vp� T�b�4֔�u{��@���Y�R@��Ci��R� �|����m�E�������k��4ghjp'C�ZGy��1cA�z
G��n֪[͔'����b
Rۚ4
0J���ī��yF�1�ݸ�$���x�m�i�:��e
����JɦylN���me<��N�ܕҐ%c�B%H�l��P�R�����v��}�W�C�HQ�zi�\��Z=�]�8@���f��/�3gBr�f�k[�[	�$��"���j����0�ަ.�B�Bc�5[߯)Al($�E��4r��t��q,� `��l�NE8�./N�L;���c�V�b�)���{�X9�A�5X@x�l!�bR��)-(VA�L�k�i� �E����s�h!@�;���/��Zu��0(�O��Cv"p�Mֹ�b��Ai��ey��Xw�:�(@bh��h��J�)��ɨ� H��ח��Wt�D�T*4A��:�G9g;�\Hf1��4���F�GvQn+s<bf��:(�H��Q�ܳQl�W*�I���ax���PGA6X�|�H����`1`p����10B$SGzH�"0��
�@�pă0�����2B'G&��*�H��0���"���31�����\��0�"##3�0�� � �����p#L1̋,��1� 3��0�`�1,#03&2�
22�*�#*ē!�,̌��I�l�i\"�'�ܐ�����x�A��$M�B��٭hp�d��eSVR��n�
5�i-�.�
Y�.pU�;x�0�M��"0�O�bP�������<�Kj����@Q�m=O��4=t4�"ua��O�n�=K&��|���t�e��HT^E/��M�v��r�a���0���[��p٢*!�%Uq�QE�l�a��r��M�=�����o�J�� ��5��P�+��q� �SH��ET�ִO<�ed�fe�ڌ�kOm�Y�[SUI�n� [xs8s����ȏ��#~^�|�����=���N����������    m�� $             !�    �           [@            ��            �  l��    �� �    	       �   8       ��  �   f����x�����۶� .� ж�n�  �  $    ^��f��  p   m��8    �  6�@�	$���հ[tڀ� � ���Wn%�� m��� �n�UV�&�-�j���ە�wm��   $m�6�� /Z-�  ����D��  8�m�M���v�I�m����c�`�d�4�Z�5��z6Ͱ�[[v6Z	   < ��^6� 	��(   �ky�-�  �m^�	$m�����m뤙�m��	�  Ht� 8 �S��@   � ���m� ��6�$m�z�  �� h   �  @j� H�p�g  �cm�q� [{m�� l 	 ��]�      �� 	t� pl m�b� C����`A ��{��KjG4䔒L��N�Ki2 �6�g[:J�Cj����v���j���8�^�\��l Ël�mpm�  �m� @ �{ﾀ   ���     mi�    	�p  -�    �m � $�  Hm� �e��χ�~/���?����V/L������i�=��n�=���+��z)�;G�/y���6n�!�O�TU���+Cx�R�\rݐJ�^Vi�E���� �7s^�f��ћx���˵�����G��G{%�6Z�Zlt˚u^�{tNBmh��9Z�qHm�z�����v�5��Rl2�Ur�m��X�j'/jl��E1ۤ��h�u�4�^��y4ܻ�n]	D.�޾�}_u]�6H�Ô�X���G�����]��C
��;�LeZ����X,{����yW�,��)a�8,CX	L��f��*���Vd�H�$Q�h   HA�s ���5��-�m��햀	6� NK�um��6��m m�` ����v�n-6 -� �  m�#�j�iW�  B�      -�|͋im ���  t� p            �`   ��    p 	 �`�C�n^� � �kE�    ?�;��`H��H�� �`  �[q� m�    �6� @6���    ���  ��   �m 6�h>@��      m�$� �   m@       ޒ�v��   8p     m���m�i��a 6� �J   �l��   �`�pp��wz� lm�` � 
�    m�6ͻ�Ā H@kn6ۤ 8�l i6m�     ۶��    YKhI�  �P  $��m�i�����'@6�b�m6�&�ٷ��V�p$    -  h H�� �   �r�&�v�VnͭͶ�i�#��a�   -� Hm��m��0 ,H�v��l Hֶ@  �d�lm�$m�6�ommm�  t kjrt���  �m�*D�� m��Ml` "��ڄҀ<I&ݰ '�i3E8�^��.�Sj�@mF��=tVQ����꾥^\t.�٤��v�h�.�6� 8���M�	["` ]���-��� ^����WmUP��.G� [l�]���O�퍀*U�ٌA��d���[���j�
��UV�Uj��X��IQ ִ�����c4�O/5�Y�e@9�m�8Ԗ]��`   ����I7m��қ�Vմ�I!"kg1m ���I�ݶ�$  6�j�8�@�l�`�$ u*t&��t-�I��$����]�6�`�h�  �koŶ�m�ӀNH �+͵l67��):vT��p ����m�t�M�T�J���KJ��` ˶�$�˻`EB�nV�6���̥�0�jp	��{v4�H\�D�ݖU��R2̽jS�[�ZУc���
�����\� /�v`q�n�ɀ�M��f��t���
btq�ݶ8s�$H  �m'@.��  6��� K)�۝� a��ւ̙�k]���|�hf��:�n9��i� �-�[R�.��   @�� ۤ�m�l   oP �       �  ,Rr�L���   ml� ����3���qn�    :ۢ�m� k 6�f� 2a  A&>z�>;������v�q  �ݭ �����h����4.�de�֤�!5!�6ى��?d�Gw�}<���P�>������D�i��8�(�.��$Q�O)�|(���8=�;Pt"gG��N�����0X�}M���U*Ҕ
�!�ДPJD#J�)��D^>��p4�)@�P4�����AlD��6ڶ���!R� � �� ��p^�����〴Z.�a0E��4�'��,-H��A���Ȃ��F�"��x��A4)@�P"�H)R�`�V�
j�: z�2�k�G� ЀF/Q��(%��ԁk�8�`'@�<8e�H�z4(ةA��5@��J�@r�� l�E�y(!�L�x�|����)�K6-��zR�M"��:�E��Њ�E}�F�8�@G��@<�<�F!�6�e�G)�\4ic��BB���y
�"5r `r��㙱8Va��j�F͸��<<��"�(�"R	"�ʢB��*�*�(���!�J;��f� U�J% �=zB����p�G;�=�!26܀ n� oP $  lt����	 � l�ړ^�є��# -r��]6/%�5䌽�<�i]u���X�Hl�ݵ���GOF�ɦ���ݓ�Ҳ��K��g�-h���I@Si��*�u/,W�v��ͳ� )��I��U)!1�tn�G4��%.�8���d-�6ۍ�[Gv�l�9�-� ���ڵ�_=橞�/�2��n�y�+	��^�]է���/"j%�G`�j��e���U�k��m���  �G�$^r�ٰx��Ô���)j�(Ջ�V�rt�bI���`�n��d��-ִ6�$��J�P�e�t��Yz\�q����7c�UʷR�5V��4[ml\����3vS��kj�<@�7[�D2�'63��ɲ�3�vw�.�9x��TpGO�����:R�T�.�L�M�6�;s��۴�	7p9K�k<Uˉ�s�GlU.aTc�7��mz�+!m�ѵ��v77��6e�c��ݞv�rd�Y�BA:mw�Ԁ��ڶe
6�ETv�]�����y[�v,�7�� ?D��G
� @�=����B8n)`	=)���eU�E�&fd��l.%�2�B(ʎ�6�#�	�O=\�+=�Y���]��?{~y�R%�a���ڡ��+�7��x�U�6ܢ=sj �;2!��t�U�M��;p��f��"f[�I8� �� �4�L�a0�k*���'r� ���!�Ə���7斎��}���v�c�QR8�+�f[����1��<�:L%�f���4�F�2zl^2ˀ�ޘ^�Y�C}O����F��D&8�N;j�Rq��0{�׮�>B4��X��(��7�ؖYKF�+��;7ɜ�����FIF��g��������]�-�(�(�vJ8�X�۳:�=T�`&#"mUn����u:Y�Ʒyۗ��h�qw�y��Yc�I�s�̺�#��֠)O�������$��d���Tw͙W%��H��e�Z�!@˜��˹�3z�˝�Hm�����S�<�Pv��=�kpZ��R,�cMJ�UYֲ�s���7�W���d��� <R��=��Qũ�Mc�h9r��@=F��(�^���CU���b��wvJW��l�샸A��TMJWױV0Z��Ew#]�I�ƓVy��=y�n���������ņ��HH��Ȇ8-KP�A�1 �lyWI���N`�]]/3$�@�&p�5����z����݊� @�,�;��q6�s]�$���j�^�����*.�X�<�F��df9��/�۽/c��hR4��U\����u>@�#H��*SqQ��l���㣄�nUamW�Os���a���p��kov�t��1^�h�I7���Ej�%+f"����V-! f�Y����L�g���K\p�{0��(�lT����ʎ]K��%��Һ3���a����1K��9�Ȏ��s���+]�9��y��,�t2�g�^���tr��qx�n���<�l�k��K�1�b���Cz�6CX�$λ#n������⪢�q�/���k1�6�^��9�}5�~D(˂��L�nNs�o�C���U�Cm$"u��V�R9Z0�U�Pz�@YjBUC���-���$����m(��;F��su^���:�Y���!c����c��&�v?:�{��5v��p7]���s�jD8ɖu�[ا��}��<���b��{6C���&⮹���jR����4���vD�ӛvl^�1EmQ�]��y$�֪�Bk�HE1�l�\H���ڗp��SC!(�,���:�����P�6it\q���VhU�
�	����)}t�
����c�����ws�Qv�$�֦fPp(�h�@�X-b��w%�/Ww)�����ڒ1������Y		V����Ň_4ǳ�,w�V�9ac���F]��UAƌU�|:�Wu�X�sd����خ��k��"L�w�����|�����O����h��f��]:���C]h���������.��K�h"���0*��E�uY!���j��M�
�Ng
28�a@��*�۱3-�mXoluA+��Y�r*{aT�6;mt�`��mt��Qr�%�.
v˝N�MT�=�o�)�A	MM��Õ��Y����2K����P$������Z]/\�����9�>>���(˗S�ﮎqt��Խk���E��.�(l�1��]χ�	o@��[VX�Mt.�!���7*X[vq-b�M\ew�k�A����-�D��N��nv��=��oK �W���wWPv��bM���'f�m���Bs���խ�tU�aܯ2�.��tR]�-��j����Q�x���5�3cfDk\ܞ�����
��l��Ō�m�Gm����ʦ�#��9!g���σ)�B�ܬ�*~,�)]��(bR���k[��S��9��������%^,��c��˂$�{�0��k,nn�P�<���\I�۷2�\7`�V�vAX����9�pZŅ�X;���l�Uy�k�p���Fe&e���=._}�@�RD�v��P���u٪7rV�ڑ��ƨ�[2�B8oy��씨�iUh!)!5o�Kt/j�Z��� �I��@�(z�9c�-���4�GbR��]��R����]/
�e�ڼ��ET=��SdN܂񌙜��m��U�},�Ё�՚,���|÷UT���7�b	�OlП	�h�C
]Vo[@�hn�7��P�"���066�c��P��6����!��-Ԧ�HCb@�Ն�+�ג!!:?����{�~��|�Ҫ��4�K1moE���6on��6�{z���4A��VZ��E�bb Zw�IE"U�%'��6E���� ?~C� ��ȿbYD<Õ��j�ttl�8 ����>��K�����?��S�3u+��uc���䪗���y�}�ϵ�6�X������	I�tK�G�Y~����R����]��������Α�&o~����~1H�j���.��ک��~�Sk��������Q;�aH:�.��������� s��C)�/�^P����?��2Վ��5@TH@x��ꮶ���e|��W�/� �Hˣ�U���ps�wjE�����V��o|�%��Q�Q@�Nl!(e�+���ۣL��s�K�PR4�Io�N�E���|�+�� ��nSe>���͌���W3���~���o����>�&'HV��%��S�n}�Q��v����
H�.�{�G8=廬{��Ü��a���s�����~��nE$q�k������`����%��8pr�F!$�pĆf!w�<:�c�ՌUl����1�/u gj���+-+�2���Yf. ���o�V��t��"ۍ8����YPjv����G�ݷ]h��6� D�A����V�	�!�;�9��1�lm���\�h5Yݏ8n�����֧
� nY��4��ٲ�Kkt��Ym���m��?~�	�{TY�W��='}wP>�m��N�����}�o�r/[���1�xԈ���9O4p
w�UU�s9y��l���[,�P�3SE-=��r&{l\�_�7�8 ��Uó��j
������Z�z�%���}������_�+2{�S٭�>fM 7��f���T��w��'B(�r��~��S�g�|��)���P��z<��E��o7��#�7{LE4�K-$XB6��հB�Qu�5W>��f���  
�	>��D�U������ r�v��ۤ�|n	����J�Z�Ox->�/�?�::��BӔ7�2fl��������ﵽ"&�%�Ըc���fxE���nrmFBC%Q�����,��pr5�6�����H�v�-=�+Xy���2��)�)8�����͏��i�:8���k�4�����i�ѽ��*����f�5���gh��w�H�&]���]�X���D�Lz�eR���@��K g,�  ͔�0�(�%0���C�#�DU�%��1�j�W؁^�h6�T|��s�5yPAե��ϲ�8.|߸�E��uY%� ��ة<P|wA�Z�S@�_L��.k�^z�B�����7�o���}gJ��ƛ.)(��z����7$���5� �������K��g��q4\����)A�C$n�mQ�{��'=�]��ylY���d;wy���fN�7�f}}5D� ��J2�<Ϥ=�ΣHվǼ�6�z����=1H�f��Y�Ϯ��t礝��גG��r9��N�$���Wc:0���M���(�%�u�v�M�W��W�V����nL�w�U�x(	Oⴞy�g��n�ѭ��G
�����.dw�jAibµF8�+Z�r[>��v�H�%j-F2>����ͻ!�(����*M:�]n�m�e�q�#�������l\�ma���'3�� ���?�{�TM������ۙ��4�:���[B�A]�Jὓ��PZ�h���mӋvÊ�z��LD3���OIFG�@o���ו���s����aN@�rbߧ�c����uM_�����=
-��C$#m˩�ÉXC3^!���:�$
H�.�ﺪ��L�b�{� �ߩ�w}r7r��ӫ��ds�W89r�dg}$�d�����}e4�Uiy:��Oh�P�)ߩ�T��EX�,�5[�vE������uB����"*�[�� �ӥ����xs����{�*hL`��#pY�˭��0�M@�w��Q��q�'u3K1J�>�s���8��W���[Tw|k�a��
�J�/bȕ^tZN!�^o��b��x�fJwps�w"���A�Уi�}��z��L���|����1t�t���%�?k-w��G>ݍ�s�'W�'_t���3�J,����)<��E!"`p�%����(����&�
 }��|�m�8����r� �R��^�	�fp 9gu��RE����"��M3wN�B[zN����a��H�Z8+ڡ���+ު�@s=]������B��ʛ)��\u��ﮗ88ocΜ�W�m�&{��Ф�Ԇ��B��6SL�������	r�zӿ=��{���� �/c��݂@�12���ꇫ����Q��^�Ž�#p�"P���gwa_�S/�����n*�^���K�~�)��߸��*�,��~��{��ܭ�ζ˿շ?3����������sf�|�oFsKޱ��z�W��ɒ��Fz��[޻Z�~O@l0�' ,���P�Ut�n/c߷[�T�)
D�_z��M�V����1�x��P� �!��m�
b+�AQ2��gq@ȌB��|���i4�bm�=����-��9*(0LL1p4�`kV{E�p|��}��* u2l�e3����M� H8h  ۶  -�  ��� [@ ���$ඤ���Z�R�55�*��z]���%�-���ڡV�b��p�j�lnVSe7���4�2S�J�����}���ZK�[�-�ڮ�
�C��� $p�Mlfiz���U!A@�I\�3���MV8a���k��+��M��6�Cm��s���(�$"J	#a��w�>��n��]�S�hV��%Zl�d�
�j�]���'mhl�U1��V��%2��<h��U����Ԑ ��N�	t�ܛf���Y:�mHsm��ia��1�*���Y@���U��J�
e00�-=�dе���r�&��_o�画`��mME&�R ���8�m��T�v���'l�mk���j�,��4�&�]buT���[l�;cx�α��U��^�z�jx/A���t���C�F$��ԡ41�TشX����*+�U] v���U/.4�r�Jvչ�NS�ci���U��υ�j��ⴏ�Yعck=$�lI4�/PvݰA�[R���+T����l���i�*e]e�f]~2��A��n��I�P�F���KT�&����$'m{BZ��j��,k^�����i�Rb�������A�Pu��)���~�{���{��?��rL��qV��C=���L�:[P��t�r�g-����&�D�n�#��fU�<���ý�&�c-8r�M�T�`����?q��<&�s�]X{]��2}���mȾ�&�g9�KC.)(�bg�o�m���V��r�����1�����3�ts�p֍��[^�ڧ�T)'��U.����}1�\���Mk� �PQ����U%���l�O� y�G��D��k�6��+^��<Q�6���Fq��(�i�v��qu�������ɦ�^����+MW �n��ٗ���۪D�zM۞F�[~)ʷ���;[w���=DV�_���RE2�m7:[W�tS^�e���c�a��$`�^��z��ӚU/��wV��׉B�'K�!�ڂB��8�Gqi�#Wb�(��{=]"�G61.�U�����@���s}��{tz��>�s���MZh���hH�&U�jn�=�a��1���*��j��'�ۺ�릓-Ȕ���?e8�zek��#۾̵��a�ϑ1w�6ggܺ��r�|�k��뿥��1����iq��b�Y��K��Pm�`���0���v�72��/������3G�К��rǘu,�s��W��޵s~��`���B�!��
_�YqIT��O%QG���f�e ګ7_7���r���T�ѺG;�����~Gv�U��.ř�)'�(<��������q���eǙ�T���"���:�i4��$e��[\9���A�{=qT�=4{޺���~�W�}��R��x��(�)�w�N��2  F��v��R_{��q8�kQ�eUs�7׺��
0F߃�Fe#~�]\ɷv�yH�I���ry�2(�-�o� m����;^��N�/;�BR�*�Q� Dt����}ur��R�0ʪ��;r��p:����Y�!b�,6eİgm�-�a�ic�r� ��Y^+b�yi�CU������uRm��R�6��l ୂ�iF´$����r櫦�.d�2�˖�6�ev����NO:������ �]���;z}F綍{�����
M���EI�(������,6�];m�:���ӵM��}��s�f���K|���9B��,S��:��w�T5�!}���./�I���� R�Wݭ�;�v��I�r�_�n���N7
�5xG�T��4�#w׳}�k��a�����Q��-n�0�.{4M�.��ip8������?rr_�?s�T>cd��UN���qx�L(�G;>_s�3�� A�.��mjY�	!�&e��"e��&j#����=ޙ�"&��w����mt�����8#,�'BjBU��}k6OS�a�T�z9���-�$����=�Wŭ���m
��v�5xv��f2�Wk�L�� ���7�V�>� ���r|a߻\m��3.�p�ܖ����u�]�V�ۘ-pw�����S�.xԙ�U�E����$��y��U,zg��d�^ʆ�]=RqK���լ�_f~��="[)ZH�^�|�W��Ju�}��UR^9�GQ�g9�#���;nU���#��Uk�Dq7R3)�s��n�k�SgTw~%C�in�R�ӂ!tm�q$) ��i���K���6�ɹw�i��{^ö� C�8[��> S�ϵ�ϻU��Ü���Kp�d�b�Ӧ�;����f�����^��aNB�4�8 ��n��a�I]J 	��I�c$!�����9	�2����0����D����^�v��8�kw���q�gԮ2Z�eUt���댲"R"�m�d&<g���8:�[�%2ة ����㹆z���юw�Wws;vǂ��c�<1�3;%U�n������X���'	�3��R���[�s�k��,l���p�)�W.Ϡ�K�*~?Uw��"�eJ���K��d�+�v��Bs$&*��ݍa�O@�y�BƟ"BX����mTҗ��U�m ����tv+�ĺ�$cv8��������s��{�)������9��e�-�VL9��!-�̅��l�av�B,�A���,�j�#�Ӡ��w	��[�׽��~:{A�a>�LC^���}��ۮ�m�d.f�m~��򿎚|�������;vWSfХ jH�5n��70��ͣN�N�3�j=
I����v�Ν��剱����T��iI�Q,S_l�S��D:�(�����یݭl�on����v>a�۝�|W� ��_�;��-!���n�n[e��B��8��o���ۯw�����[s#7�R{��0ѐ�u|���͇���s��s]��.%w�����^�#��lv���%@�%�=�5�NG+ي���&OC��J��$�}�uW��m)y�U� ����tWI�9D�Y�eWH�#W��/Zʦ4f���H�Z��RF�ƹX��e+��b9)�W��Uy�����ҙw��pW}1Ϥ���P}�5>�� D�g��֪�������Mbrg���P�pݡ�5���ݻC��?�/�竧G�kG��_�ַ2�k4q5���Z��9ó�8M����Rv�S���*�UQD�(�E��h;�Duj�أud��+o%^p�\��%񪗔*�Ԯ�����*��J� ��"e����i�\��f6y�v�4�m�T.�,%�V��J�b��AD"x+(���㢲ʨWQ�d�
6V�NY�kFM�d�����He�����5W��b��^�Ɇ"�j�`ݕyc�,�K
|@0���O�B�`�R�,���F��-J ��R�V�"�V+m1�`h���oB�ښK���v����J{��� �9�S�*"�' �D�$���H� ���"���I�&����(����m��cM9��j�
Ex0�	d{�#�6�����D��hg(U�Ugj1J�%T���ܾNs��,(@,���� X�z�l�i1)�5�X������s��Wj�?:ڡ�Т:	�]#읕��˴{����LG���E5"J����]�T^xv��{R� �u[E������2jZ!����;�M��u�oӦ�ڃ��ܪ햋(�7^n3M_q߇lP���c��uB���E��)H�(Mu�w]h����8k�j�/�U3}���F�k{��X��S��hpã�pu���;p��  ��٪cýM8�K;%:�*�q�H�c�~���N��b	��.#���e�e��ͷ�l��w�_�!��!r�9$G��}u���Hp��	�/�T������F��{��fm�m�Sd���^i���L�8�a*�"U�"9 *W���q��K_��T�-O]UkE�눤�a"In�ΩV�:�ʪY~���"�h��Q]P2S-	�3����$��HĐK vz�환fm[E�[/������z�&��F`�i���KY��1B�-��{~�vy�< 1�HS,�t*�p<f�r����P+�u��s�/Q:7��̲���,�Թ]�չ�ܻml-�I��1���q�k�T!����@�&�f�KEc.���!��W�UX�i:�|9�o�'8 �<�.��6<�h��^睊�LS��j�����[8�*I#T�zH�Z�X�ΧÜ�n����i��8E�!�9yOi�����oÜ3��?����.�>Ҭͪ���6���su9���/��`Z�Ô5i7kG9�=lV�J��_�E�Y'���pA+�{��p���T�t��� ��pY�vn�_/��}����-:����"ٷ���*��"P]�wK���(Rp5!�τ�~̠�[*|�UL��]#���$��ɚ��]����Q,h�u�]����ZJ')HY[q�z�_�Pݩf:�jh�Y����Wk�ޛ����v����8�f#v�4G��˪Ű��U{�{�<Q�[iz�0_c��ۺ�,ծ���Gi+k�\�s�0ёGuk�Y~4���D��O�rzNʽ;a)"9*��}3*�@^v]��}�kZ���\T��E�{Jr58�E@�`u�[�)�;-� ��[���FX�J��.p�۩�$�G�;
.H�4�����U���UƱ!#����[̬{�˿mR�WM��]A�ܻ�޺q3��)g*w�s�=�Q؜H�����ly�m�n�Z�j��j�n�Y��̴���	����A �������4� �B�1��r��[��UI_Wrň�����OSL�R��D^I;�F�`.R��_m��mI2����w-Ȋ�N���},4�u��c)���o��9ْ�=uV�yTW�B�����~ͪ��A�����럫3�Ȋ���_�w5R�fa�U�'`�W��֍������:m��a�tA�X��pr�!��9:�����t���4쩶�yzvxͨqٷ��y�ň'L`૧*Pqq�Wn�
�W����r�m�lZ3�FX�������<�g9�R�C�I&.��UQF�O��kps���{U�a��= �^o�T0���V���3�N�O���qĕ�ob�1eW����m�;�9���]�P}Q�[iC`������.��c�K��a�"S+:���ݪ�n��{�W��+���o�3�k,n|^�n�\)0���e0����o<�@������^�R4�\	�I&Iv�|�y���7�(�����S�̯'�&�E�Z���n��/�e�e����N���l.ȑ���}wA�Y6�Ƌ��U����1Ḣ���o� $�S0���D1�9�n5�w�ͳ��o>���@�m�gfV�eB�hY�G��o�<��E�������#����|����y-�z7�����=�"V�M���N������h��$�	��5 ,P ��X"�(($�	f����qۭ�5��]ҫ�m)�h��i�ڒ^[o�D���1�ʪ�E��3+̅͘���?)��v�=v���%gHp��� /	M5�(Z���.b*�D�.B�[e���g�9���}�v����熣ऒIj�~����6�y�����U�;�fɔ�q�iwު�ꪧ-����n�m�{���r ��^ȗ��wM�kDȶ��1� +ޮ��{́�B�JP���얆m�%�Rkn�e|��'p��Y��ˣ�3��fg:]v�.B	6]t2#�뿞�����N���,Wt꧎Xj��8\�K<����M_�e��E�c�A#�$ʕz��VSKb�����B��m�SM��秽㙗�Kr8R�)���OaD7j�}U�o:����={��2����녑9fg�g�����¨�+2�30k"���M%^�$����ז���p����6�,��EhD�sݥs�p�kJ�i��@1�y)l<l P���!��0�1��g0@�
4�#�@�0�	1�(U���M/K�A�K�.��@a3,���"h�-�Ȓ�?�U�5tr�W;�.B�$�'����>"��=m�` 8<�m� ��  ��  ܲ���l j@��"���2�F��Sʪն�f�r�T��;7v��8n�ù�4�u�cg�c�C��˚\7UK'�j�����=`贡=)(��HpYj�@��k�H%--��'�5U>S4ʣ=��t�v�֨5�4�o%u���t%6� p�e�Ĳ��C�/-�-�|���+k�B���%Q!JKju����o{� ��]�m���"�(�RI"��uZ��V�B��4� Nn�ki   p'G�'+U��2K��ej�.�Ij��i�.��`Yv�K�)��Tધ���������$xi�h
�	8CU�ٶ��Bj��ҧ1����mUʷR�56�څ�[�ː׭�l��H��FU�p��cP���J�n6���b`��Cu�s�mF{8���S�V��;t�S�!���8n�'����V)�َ��r�'*'a��m,a��`tk�.`vI���:�W.�-��Յ�䃋�-b�[]�]����'@ ܶ�
P6�7i�4�UH�l�S����|(����ڨ�P (�; �[A��b��)�SiB墁�=�߷�&��$
���k�g���1"э̵�)W��h�bqٍ��5C�����w;�:�V��ԙCkqw5��A����1�+ad��h��e![��Zjh\��m^mrl������D�M�dWlK+���S 6�[X8��J!�١�p��]������}^���W���{�.ڑ]�oSq�eUu��>�e���r焁�(�c[����۪K<��ݤ�����&\*�X}�λ��*%�R�6��9����p��If)]�}�V%k��]ݴC^`��hn0�b�T���vv��.m� ���jDE���K��F�<��[��T�+�o{CUy%�J��W{�mIt4�NY'Ƃ�૱)mt#^b������o5jܺ/è�Q���k}^�gT��I���ݡޞ��3�V���vL����]������(4��+6R���˻�E��UQh��፷a��.6�#+��,n�ӎ�c��N�
���J�ۯ[{U4��w'�l�$N���m���.�<�@ߧn��Ұ��2�^oU2��f��uہ�ȨD���2A����ϻ[�s��{�D����8=���N$�0�a��ߓ�ʹ!�ޱg��> o}�aWH�_.��8��y]d��f*�g�x�7~�q�7�r�j��a���ٸ��p�}V��MBe6��k�!R}Y&B]����]p�[z�8Ձq,`fk��cW�*\��C�O{��n���Q5���ϣ��29��[�Ḝ���C"�N��1ɉ�>��f�N�D���r�B�_r�G#������C�PI����<ˀ��T0�a�!�Lq�B��n;�U�{.[���{Vj�p�x"�I0Ү@�lC��b�!@��}�~���#�eY�!�h�7 vx�N��`(P�؅�,0�
�Z����k�����V�C#\��ׯ.�&h�wD�.[���>���5�J�Ù�i���,�r�g�(�b�0��ٙ��]Ԓ����r����%��r�^K��ͼ��O!��ߪ��؃�r}�K�B��~�qܓp�}����v_�D\)�x0�l��G����w�9G���x��p/�U���}2�r�	y����C#�z��q�Oe�r�ῷf�n7g��Q�.5�Btt(���!V���9da�%�>�g���2s��.�.9��!�![|�g#s��L=������M��D�~�V��MF��	3��Q�.5�Y�乨<繏!��\�l�D�ϗ�u�KfH*ͥl.$��U��*;;]��4���cME/D�u�E�D���[;��� �t&Km�ε�8{7������lm���\2Я�Ak�\&�+^�v����pA�e@x�+���ܜ-��y��Qm��}��\*��^�f9u�^9��/�V��F����Gp�N�,t�HC��3�Ş
<d;�S�̄�Q�.j�m��5
��wx���NN.��� � B���g�ܯ$3.�4r:�"}�-�\���5.z�9Dg���"��|��@��&�8�'�f��}V~���/�V�!q��b�,�"�6�|��<�>�ZpA$��97�w��7��e��CQ��;�NaG��Ɋ<x�̔�D��A{
Vݹh��^����&B�n%\�����,��9��d�S"du�و:����9��5P����~j�*T��C�=﷎�yfŞ\���e�W7��܉��=Vj��y�G��yw�Y���cH���\23!�,�x��LQ�ʈ]a|F�"}��d2���������#O<���a�\�"���H�B�< 3�&G�ݛ�ḟ��B�\u�Y����?^��D��4Æ�0�y��x�(�%��9�CO<{I�<x�w�"�I�}�柼�M�_�38�H0���뫇�k&�Յ&^{_����?O�d�P���Vj.�srg%��O�yCQ��Q�jn���˻��ḗ��S¨�7�_*�㑸��w��.[����&�fT��u��y����LM�p��ܳP���pd���3׼��7�խ{P{���"�!�����E"76ŹrJ���w�{���Ḟ˖�.2}�5���PO~�v���c�\k�����7%��#O޻��,�3�D��yI��.�.9���n;�����S���1��=\�zvx�6r�me�0+����N��1Ɏy��:8j7�e���d
��j9��p���'0�<��t{�Yn�<ED�L\���r��D�.[���wLQ�O,�!�Jv��k��,�x��j9D�{�wÏh5_�en�Q�]��.9�#�������U��l�I;�nB�\u�Y����Zy�������DP�CU�{�)�<���r��ޭ�uz.Ufi�7�}�[�����iq�\~�,�w��\�'fDÝ��,��Q�ڼcdpE�;�M �x�+�]neW���זQ'�}-7P���f���O����6ś�@�>���9D"�v;D��f*�g�����f�n�����n�ģ�FO�z��\�,����&�-����"~�����9#y�Y�����Ն�yDC��g�E����K�Fd5�#�N�F��g ީ�{]���ᑬ�y����tg��o����mH�dNFꋯ��㑹�Nr��p�Oe�r��j�D*�F���*�RU}q�*���������X�C���.���V�����{�"p2�b@bDv�[գN���M���cn�9���8���Tgv|m�����X���^s�c����kn$�����nݦ�ItVW�Ֆi��u�s�s����k����;^l�iR����Q�#���$�������B9���EΦ>������|���ל�
�
"�H�����7�٨C��X��r��m9�[Q>�z)��jJ�G��X� �[��q_������FB�_��!��ռ�L�w���yUW���r�I�(��~��&�q�����*|�PԐ4��澖nP������%]hdw
��z�P�*��[��>�0�T7M�S����k��m陴\k�%ճŝ�L�����Z�.��}a�ٸ�N祚�T+�U�����{c�j'O��Iz��֝¢r>�Vj!�6���]T|q{��hd*B��dC��͜���'F��$ˑ#F��7�e`�G\妧�n�]��}��x��O�̆#@<Q�޷��2��v��p��� N�D�S B�Y9_�L�\h#��]�
�E�uf�_��$�F��;�G'�};�ՙ᥺� �hCS�"�h�G-�띓�o�f@*5�Ձ����YQ�5��a��R֓��%#�k���H��m.\2'������K��n��6��)��U�,�k��>
"�u�d*��!BCһ�'ڬh��z�<:;��JTTU!N�1�m�n���So�.ׂ��b՘P�&$��a�u�A��خ(k,dd �A�j�w�t7��:C�6������#+�m�B�&č"�(=J��&@Bv��$`k���10 �H �Fq�"#�� � ��c�R\�"��0�0p�qRL	�2��1 �`���̶�6��.m���[�3%�v�Wqf�ӭ�z�N��Z�V��-���։�06��D�S�t��֑D�iT��P�|ɚ�U�ћ]k�r ����!�״�7mW!�"�w��5 ��Y�
�/�ա�~[��i�Q���y��er�G�oш@�xX
��o�>�.CP�wV[^n�FG�}�n횁y\v:h�؅Q��rw<>��&��OӌF���ϣ��q+�nB��,ȅ��#�B1���q�C��|��>Y�oň@��LG���ָ�fV�Q�N���T_ʳ�՚��Q ���G����}c�)�#nJwD;���»ڵ�!Q�ܱ�5� lz����/��ܷШ{�KƓ�:y�Y�E�B<[l#�D<�|�(�-��B D}�/�k���}�ܝ���7G=�E�Jgʃ�@\��`!w�>
"���|��qw�VjP��-�GW��w����̇'�?}��������"�� �#���x>���W̍@>�Y����hc��-rHTk���"�|�(����Ҋ%B���8_�V�B���]����o�nB�j;�>Q "��Rx3!��@4�<���P����g}���`�ՙ �W;VF�PE۰ ,����uYRY&@U��6�{+��j��GV��C����z����Co,������YO0�Ba�d+�}��gU��v[��vu��VS��S��IFm ��UM�D�2d��\�B�y���.��a�΋Fx]THR�WMtJ+��J�:�K�(����j���܅@7ܳ"
~,a�徲x�"��Ѝ�r�Ho�@i2��6& �"H�k�� <��D @���I�T�F�U���hd*{�L��χ�"~׭�5@�z���%��;�=����@n�eC�߮�p�{���q�b�9����� Q��������q;�[�j[�Y�
�o�2��J"�Dӛ������v���^3�n�ǦOS̷�߈T�e� �j�-|M��~��<�_,� ��N$j*x!oɛ�G�a�v�}��9�-5B�w�n� _�&u_gU��^cm3C���(��(�;*d~ϯQ.�z�DU (���y������!/u�^]�ei5��܅D7ܳ _р6��r�_<���=�M�NW=�Y��Y�~�=3�U��T{�Zj����%$�|���o�;F[���bH10B#M5فc��\�w\���#'� (�b���DB9��	�(��1y��\��T ��y����"Kʷ!P��dB���ZT(ꌇ�3ꇍ�uy��n'ﾷP�B��"(gM�+�x����7VAv��9�C�G��FUr�G����՚�T7~��q��ҡ���)�{�|�Y� hhޘ�QD�Y�(��<� �!�����a���!�8BIH^����yv+3`ZR�m����]f��(�M���w!��yZT2'9�u@+U��:�X�W~LG��;ZI�+�����7�<��E�f�����T���s�<�١eJ�D ��� 
�s�k���2=��bn�@��~EY�J g݋�'	RJ@��	Q��ơ�7�א�*j�Z��=E���#����R* Y��MCQ$�z܅�7�Y�R�d9���t�!�g7�mؐ��0ۅ��x�+	�x�D�M�cq�����w�[�n���"T	
��hd*r�������{�Ԏ'!ug��@�ĀT�V���Sp��I�Q���}�� ��������xj\���2F���D��܎Cpg�̀T>�������b��3G��r���W��h� W���hQ<�iF����8س+I�{���nC"\�VjP��X
��I��&�$�F~��,�61U���bܴvc�Ԁ�V<����Nz����Ba�a����1�>�ߞ�����W(����WI\�`��-m�u����sf 36����Ё��+�ZἮa�w%��\�`������K1�W�����z���z-�F�j�v&�ڮ�D�xc��/ۦ�
ߪ��Tw�Y����^�����½ةJ;�#�Ł�D`Q���V���v 11�,ƌf0"[����C�$k�ՙO22.F�r��A�`2���^.��^պ�CPy�Vj!P��,�F��<$M9\�0����"� ��(*P���G���Q�O���O����K��d��fD�n}�@�n:�k��j5[�:����˝���cW%�h�n���9�'@����sq��RDhY��c|��G���(ٳ����D�y��$�����fl��G��_h�Cှn���kFg��|�� B�������i�R:��x}�~.˻��Iğ�nC"�9�Y�@�o?KCP���iQȜ�<�\�R�����w>�jP����G�妡��ܷ!�Pr$�&���Uz��JOw�I�s���IϹ�U�E���"�(�p1��Ϯױ1��m�m�lƴ�nl"�KX��U��<%9�����:8M��ۑ���ڳh���/�`d*>�_��ʅޒ���{��I���I�zY�����X
���ӹ�7���2����Y��� E�/�pAق�XE�%Yb �o��0�"�w(� ��4�Ho&��*���Ty�Zj�>����|�@G��G_B1&� ,��ip�=�-�5 ߰�Z�.�U�����{h���p���f�F�M�ÈeW;L���D�'�@��C"v�Y���.��`B<YlQ�<����M�NW,�H=��Rjz.B��hd*?��MCQ'������9#�d ��� �Tk]�����ϵn�>�̀T9�T5�[��\�d����(���d2!ϲ̊.o�z�k%�a�\yyP��2��4���޳�p�$N���!oɏr�g�f�
"�̚��`G�+�R�SWh��n�l`��xD��|�֝JM_e���ֽis$��r�CP
��d�Iu�0Ѹ��HȬ��ȴj��a�&�q��i�ٸ�����P��d~)2�!��K���^M�Ty�j|庆����ĸ����GG��ڒ�(�4@^��"[� �����@���!��3A$��Y@��Y��7�j��T~�,���Ν�PN�!L��ʂ����.d^�j]�h��'ЩD!����ef�<�6�I�.P�U�1�8�Jv���{����y�JS ��E1T�
��IK�``!�%�Ф*��@�Л ��	J�Q��Er�C�S{��-�Җ�%1!G��pA!�%`����at�-qQCA��Z:�0n�
E9m:	�(��#fA�;H��I�$R���nI	�)  ��� �` -�  ��6�m 8l��E�$�a�Sm�\ Z�I��e�euY�����d��9�u�;�&͌mbqôV�r�Yq�fe�H���9#t�;�@s�����^X�ʺ�b��@CUIŲ��*<��z�:������NҪW��6ۍ�[գ�7m��H#m��)�bVu�u���=q��Z�R�3��}��Q�ӂ�y�!.Bʒ�L�)�J��10
���Yhm�	�[m��  mp�,b�ٰ������%���[Kt8ݰ�'Ce� �UFE���
eJ����hZ55 a����7,���CCI���L�Լ�V�V��@s��.�@��wI�kYe�Bhc6���W.��(ؠqA�Yu�j��1n�*�����k�� ���M���hY�m����8�йG+J��TS��;e�v֕�� �wmVSw^,��k4Υ�s2�`&U�j�܍�]]�TK�=,"��j�f�(�j������8ۀ�㇭���eUe̫��B#�hD��[E�K��:�x�i�"R��{�r�S�ьN�u�Gh�6�	�:�afX�䌲�C7^D����J�Ǹ޻�c��q�Z��m�C�d�[�z9Q8�c'\ة�6�3hj݀�y�r�[�]e��t�z:Y��n����A�|q�Wt�׎�ѹ��GV 3t�7l�A8A
4�1��*�T�d ����\p��]���r��.��=��	���=v}R����G����5w��2��f@*���X(;�C#�a^j���w��nz������C�iq	�'�(�y��9T�<[���Y���}LQ #ӓK m��1�DB�����F�u�"�$��"\/�U��J�y�MCQ&��!��Ϯ�$�￴����f� Y�s�y�F��6�a9!�ї�4d=��d�i!�7�oTj��� 
���7�+y?z�חe�V¦�ș]�D5�x	Q D�$R��ҧ�w;�@>�Y�P�G�q�!���m�NW0��	�h�z���/��_MF��=f����!�1��|\�2�Y����E�����a�P�}�u@;�/�D �y��\��T �\g��|E>P'��u
�w�Y�
��a`d*>�O���e��-�h��M�V�JW�\�M�9�'`JOu�!xlB Q�L�_  M�6E��4b�J�d" �ш@
�B���ҡ�7�[�h�W�{'��3&w��n��`d*=�m5?� ��j团��y�v�@�b!~��f	 ,�c��Pț�-�5����Y����V�{���y����i�ܕ�DY���_kN�Py�V�����Zz�q��ґ9>~=-v�
fkc,v{����k3���-42�3�;'q|N�d�.7�j��T~�,�=�5AT	8Iۭh�|���w�q�ĆIB�,�2���C-�9�P�N}�uD7�d��d��ҥ��Zp���Zj��]�
�l�$g��� |<��{b0���zJ��{��P�}��5 �W>�!�G]��ZI�f�`��8�W�ݯr�y�_G�׵5�b#+�B$��D��Vjn-����-�M����C"3���в ״�
��a$���ڲw�߃�u%�Uk����2�Y�Vp�и_r��G�妡�7M���4����1���3#n
 ] �=���D{��ýo�b@ b*�*�Q���K�?z뗗e�V�MC�"_﵎B��Y�=���,�>?m>E
��/#"i��G��� �[��͞Q�9��"�T�yO�B f�5!��@�����$5�v�CRE�p�"�T.Dထe!��$	�w=�%��UmYc[�m�K�x'i�\V��aojڝ��H�%Wq�P��:�t��'g�V���9iS�{.oK Ӻ=/,E��G��Y���{t�������7gFc/]uh�l;��I:K�oj�������%��p۩����Ь�Uk7V]}��<&9�|��5�:;���p��������P#� B�Dh�4�p",�o��w>�<���f�
��2�k�/���������NL�j���۠�۳p
������P�rҡ�7�[�j'����\̘j���B�}V�Qq�i�j&�v�*'� ���ܳ�
�~'�.�0�4�Q��ҡ�$�9n���af@*�U���lD�����J�㇧˖9���g�v��G�s:7\l�ߝ�{nIlf�b�.�.��ȓ�W����s� V[��5>�=i�.��M�$2J���⵬#�9U_�����l�ɐV7��3&����ae�Ќ&�!�Wݒ�K��gnJ���J�	d��h�۵����\]�v���a$���}��@z����`x����Lǈ��G
h������Qc-�!�i�fF�mir�L��9���@�,�IM%@R�D��N���3��FY�#h���E�f�0�n]iucE�jIT���f����p��ͳ�<f�h�,�yh3�h��� �q�kLF?]���y�ii�+�J}�7x��8���F�۪ӭ_���]���%KZ���"��]��Aig�ĉv�Դ�MD�S&bg+�����Ё����/u��vG�,��{�n*6�C�ڭo� g�_�E�y'	/��w}�rl�� �KDbia��0�|�.3�jt~4���_�SL�$�ާ���3n_##K��r��[������܂��(+�q0n�&،�(ZY��-/�rM�У�z�Ad�(��s1(���^��¿�+����횴!Tc�����ՌU��<v{Q���\aǟf��g��27<�lT�n0�󿲷�;���kb�y�-Ul��q�@\�BtL����5l��`ĺ!D
B��e���c�2F��e�B��&�x�G��y���mn�D@�n ���ˌC2� �c�٤ۺ{�ט3�1���|�[�Po�פ�A�o�@M�f.�CW�^����[���(�0̻� +���[$w�S��8��������ϗq�q�ȉ��o,�[�����L�AF[�gV�f� � B9	��~3b�&���u���wܗ!�v�k���#HrUg�g1�fؐi݌Z9���d���]�+�GX��ܙ�R���}�Y߻$�������j&���t�eJnۄ�S1Z65N��RV��q�[p�WkWR�I�Q2�u�X�(s��R��p]�9��-/�7�DۑrM�n(�%fW�mO;6έ>��s�w������O��-�3����urm�{�ʄ7�L�$�nN��6w?e�7�#$��T>�%�
՛]�w��P�D�h������*��Z2J�*����	X-�@K�p
��9HaW��x�B58��C.�E�b���D�F�]�A��o�͉)b�Ӡ�M�(���&� A�胎 0E�X2�)�9&����2��$�9���C[o�	���
�}��4���uF�f�/2�Z�ͼ����D�tO4�����j��G`4�@����-��ۚ��������\�w�f��<�D�%U����\�1�����%�L���88{6K�*�SN�!��|�u6�N���fV���� ��&@�g�Hr�<��S&U�&�!�]͞��Xg�ĉz䚯�e�Lj�'}&�TƬ����72$ߌ�`�����d��#����*׼ �<��Y�E}�O��~����pts��/>a�c��a��\^)�4��g��N��t�6m�1��ڎ2�;�Wc�l��,/֎%�@�s�C�ĉ]ȵn�Le��a�	TNjf+/�rV��2�1��f&�o����x�@,.���z���6w7� |/���((��3�ܟ�}=����UP��ҕ�J��z�p=��B�WCb�-sLH�n�[��/���;{�ʙ��pk�2Ɖs�W#�.�e,�p1F8���mh5��e�����qM��h�B^)�HlXw.�����'�BHI����뻷6\��6�^����^��V졺vc)�o�UZK&�=������� �{�$�Ɏ��W�>±��R,�{�<��W�pp_աX����P��j-�ܒ�z��d�ɓ�����+�7�(�8 ���U��9){]˿�B#��in�a0���w�'��H��Ud�&NU3=mI睡F��s0��LÛ�{?�0�I�����6 ���9���y�īQ�u�_NԌ&�,�_��V0�s�������Ӛ�G��cT�}%��3����7/3���R�'MG
0`k�'��*
���}�7����1���}uX��ˇ�͈��R6��7$TR�S*�U��q�z��c���i:���Sb9�ɮ�89���8=�|SiIwK}j=�?i�@���<��ن���7��N��ϞM�z���&���;�V=PDЪ�{�	�ny�k�"	��,�k���y�t]�Ή*����LIW
���K~o޾������e��������s��=&��M��s�_��8/s��?P,��ʼ�%*�A�kd�ʶ_aeH�N�W�n�5�/�O�⌻�E��4���2ń���e@�h���dAĒRCe��EUS4OG�r�7�� s�  �{������-�㒇��2e*]!�Z�
�(�����IA'P-�Ɯ�j@�"ics�A�UX�*i{`ʾ����e��q%�]3�+�����Z���M[ ��dod�cu]��]5��M��-VwT��3�c�R��,�&��0��;���n{*k���;����;*��%����8,���*@�LJ$�*��c��%J$���F�F	�vĉ�"f	/Pq��.{ꪢ��fA\tC'e݅m�'��;8�"�H�؋8x��)���,�g]�u����h�E���emM�
�]m��:�αq;�nL��X�Ig�C��V\\ؽ%�˗p���K�2˄�Lb�T����dzX��+V�V��-�ȹ(��/�Y�|��9��;M�7���
m�h���MU��u�qw�O�:��6it��b}�zSiIuW��c�=N�v�=o�$�<�Ɇ���-,���W�{/��_ ���i�c-��b�KMD�@K�v��Ͳ[�ⱺ���ϋ=�M�}�����gh��cQ��>=���� \d$ ��( !�=������@ <��o�������SJS�o��o��S�\�������`�9��M�w�c��N�d�
�[�f8h��b����������3w�Q�4�9�qs�:y��#;j��!("-�㒇u����s�+l�y��J5��~�~��5H>�� ���H�rY;�ɬ_�� ��C7z��{S�r ߵ�s�Yd�.�|rÐV�%~ ���G-|��R�dզN�[�&�,������po�C�Z<z��_��7����&(�K�ثh�<��6��Y���
iИ��6MZ��Nm�;����F���x��OS����^���m��7$]�w���s��У�ͯcX�)���b������v�M}U�S�D~����@�=��-��Ғ&꯬d[��o�N8�xH8�%I��D���)"rF���������Y�L���W%k˵c*�s��q��#��ɓ]�F�f�Z�=��ܕxB�\�+�C�~�2o���;���x`,��fv�v�ػ���j"BU0�T}�]6J�g��0�!ډPj,��|�JH&�&�P&F��%����u��I�o�+�4�9�(QF�G�(�1x��42 i�TGXh0��`�n�M��lB�0�oF�.؝Z�*��! �M�L�c0� ��f	t�/0��+h��@DM0MCD4�Q1E�D�Q]t�GntkY��''���*��IU)`�L������0$m�` 8<m� ݰ m   u���`� �[R �A"Ce�M�'n���]�×M��v1l@t�+d,7U��,E4F���& 6�x�I�ܚ�f�c��X�X*��e�%Bo[P�������� s�c3O/6��D�Q�v�ʣ9���'�Zc%G.����
�f�P�UZ���U��85������#���a�{ޞ�O��ġT��z�����R���v�f��V�*�&�*�vDLs�H"P@�-+Z�k�bԬ�O
A��e�I��m$  �$c�I,0���:�ֶ���v��Ͷ888 9n�[I�m�wc �h�m�&�	h��ۜ4jkN��;t�����۶��m�mh�*�[�@���hn��vMOl���������:����e�Ytu��nz�%���F�W-�W����w�x[1�T��v���]XxE����������8F:�AՊ;���Ut�탗��'�7�(K,qJL�0'Z-OW���ۢ�e���3p�*�[a�� j C$��X��r�3����yX6�t�V�����H�4��,䗓���
h1\@ ���E�,����1��qG`��{�&����JUcm�l�K[6�h���o6j�ҩ!a�=���^9k�C��������b�y�3]%gNNZ��f�P%.BSU���+��s�C��v��-��u��3Z�lq<Ƶ���ul6��s�q����b�yha-����sٶ�Z���Q���W��˪�,\Y��D��h-4��ӭLn���t�>Ox�9Wg�3��pm<Ϥ=]kyy�n#$�w���ԯd�꼮�?u�}pFK�ַ{&�jcd�W���^ ��	�!L5�m�g��Ml�͒�e��n"5~�������]�&���+���~o�� � ���~���{{�q%�#.�6�s3�z�n$FK�6}W��(l�����;�$u�=��{���Q�V!�s�8A���.������l3�ε�O�:�ֲ�v�&iQ}$հ���G�7U�p���8�v0���%��v�u��1�{_�۾b&�S*d�+j�-���U����/�ECc*�����ia���w~���ME`�_���ۢ��������(_�CZ�g���qU��f��)�-_^�� ש}K^�׋����xy"<�T��x��=��u1r0d� �>�z�^����L��7�aR)J����V������������Cm|6Q�Սk�V���)���{���q<�@�����Aݗ5����k�
>���?~���� �8x8.����A"�,3U?g�>�g�l��sd��z����*(�N0� i�4�գu2Bga��HK�-c�L8����F��5����]27��fP�3h0R�2b��J�lm�!*+Y��i��"���y'��I7�#�d5yÍ|89]���y�:Z�)wZ�����M��y����]��/���00	Ɛ0I�Ҏ�qI!8���$����%���)UBڨ1�,v�.�`"��t�hZ���OFn��1�ޕ�K��H�a��z�Y�;�嫡�80�</�^ms#Oc�q�]���ebaj�gAe-E��*j�#g�C�z}q�j��L���rNr�Ü���P�n@f���"7r�0�B�uZ8 ���99'>_���5��-��s��{�JH��ߺ$0|��ⷒi��p �.ɇ�ʅP'<���Q ��sM*��>�j�A�ʂ6�{�5�d
�؈���p%}L�T,���)�R��V��v�!��N.���D�_;�vYKz������&Ņ�B& �E��)�-f7�>��P���ַ��ɷ�>�.ʼ�N~��A A��ן0  s��Ϗ��6MyX~qB�J����f8{���ϩ��tvd*IXu�1�k��Η�Ǽa�r��G:�7�����zh���(�F�b'f���Щ`x8z�r\n���n/R	7k�˲��:v(}���IJ9���<�5�;Z���s�E7��ڽs�_���UA ��j���^��i�"!K��nz�M�m�WD%�����Bk1x�ۓۻI7�%�S��ڄ֦}��:��8_��@�m���WM�����Yx�)Wd��.��_�|�<���}��q�0FI1��x��Z��U�}�?t��R$��W~�����,�I����&�|�TU�^���X���Z�5����<aJ������Q�,~�*#Ukd�q�_�&�����5���p�0Y�Ҹ�����!ħ�`p�S���.�`��� "�}!���=�<���c�~lV�^�QC/���~� ��Q�$�^����2�r�}���NױC^l��X~fD�J��WjJa�����k��ܕ3%ff�v�~^o�Ԝ����F�<Q�7Gt�øx0�5��8p�g����
�i[��B9VP����r��\jV�,k\-ሷ	`QC�x�k�篑임 �j�6��W.��d7%�6خ��з[26�'��R�;B���v鞵sIt��	{(�UP�R�2˄?�
	5�r�o�ٺn\�vv��姰.n���XJN0؍�����f��L��ײ�E��Q�:�1���w$�/hS^z���$���U�D�m|�����DB4=�&��*>�����ɹ��
脨�_��yj�K��%��!B�P��-P �T�0�-�Ӛۮ��QF��-����C�~����@�j
8����	�\d�DVAb�Q"��ڟ?�߳�!� �s���\�2�|���d�;��m�[���K5Ob�%6��*�]�Ծ��g�7{�F7{N�xL=L�UE�;�w�^I}a��l4�Dg ��8x|�.\���:H��8����HV��u�]a�4Y�b��"���Ό��.q�#���/��$�L��o��V�g��;HA�.�/|���R�41+�nn�Ѯh=
B���*� PY@�tD��w�8E Q@��c��)w)209Uy����&�V1�.!�SL(C<��5��N��u�-"�)����h�*��)�31�\j$�! ���%���fY]�j�)ז��nc엷G1I�9����ƄB���i��"�/Tt6�!?���9߷|����U��p	~���oG�-� ������VEvOb��X�>�"R#GZ���U�xg~�9ɾg������ˣ�5uټ���3�+;�}�hz�j�U�Ll���!K���q�lF�U����is� ���GZ�\	S8ꥐ���9IS�g�'j�a��x�l�FLֿ2�J֫����5�wY����S�Ms�3��pp�K��5��Ȉ�7�3������ߪ�1k!�%�Ki�\ ��)���b��a���k
�J���6��Oڌ��Lܧ�Hd1H,��~�����g�ќM�/<����2֯ۼ��l3Z��W�!��&:Z�/pV���w!o��m"J�y�k5۪�-��{hY�<$���I�����a�*�������������t�����8{<�{��]�g��ߧ�Vtu��n�5XPL���GN���4��9�ݧg�&�;�K�}��nK���X�j&6���R����Z�r�����x����nS]TX�0�3e�d-`a�8���
Ӌ�qR��w�T��3Q"j���7ݩ�L��C����_�_ &P���(�p֍앬3_;���Aw��*FcT�;!��(ia}ō�Q�3G`M� ��l�ٻw�ڮ�{�����5u��멬���f��0)��Fb6qx�w����~�HM�_ǲT̕y�/���}��C��HB ¥H@XF�!"��"N�����_��������/���A�㎅_�f��89�9��(�F�v1����9�Gs��c�=g$��ϭ�e�� ���%,��ً�"���@�ڐƺ�T!k�l�p����
TyPR\u��W�4�ׯ>�[����!"H��FJ>��������bN�9��{S/�����z�C��y��]���@^�:��9�s���5i��1���@�q�/���#�ˣ_�J�;5�֐�h²f3ؔͪ4�Ȓ��ڶ�X\|%H={ޝ������̺�ї;Y!-��I\9��
�3��ڨl��{��a�2�Tqt�ѕ�V䆵>�8  ��&�Q"j��窱�#���n<~,�C���NU4/�$7i�^������~�9��ղ��z��f5k~l�<0���ܘ:��'	@���V�q���Bz�Ğ^��*9��rQ�ѡ9�}�Լlo��Fb4q{T��uZ�(n�3_F(���*��a}{%����6��`��A$uU�l�@j�C]ȥ���A�FI@�Xf��ܐ֫��=�Ns�����dII[D�Yv:v�9���:Y��'F3X��I��[�Zj�Q1�߾^���w`y�e�D.1�A�=�t:y�ٹ�A�]ces�+,%��^��\̤Ad�e5���؎�&�̤1�Ne���;;
\�zx��z��n�2[�-��x�{%k���טd���&B�n��!�L��W`���@��y�5�?���u���z�C��ſK�;ʮ�Nށ�/�:RCu?	m�(��s/j��3}u��6[L���X<���t�w�v��ܭ��F��$IO%��X� Ϡd�Lz��,�"J�W��7���i����Wr��"�~�Z����(�?�*mg�3�˞�>Y����mU,�T�mO?CL�����fHk=��f��۾���(je4���H2�}<��h&]��6ݕTъu�O~����P��N�>�wA���Tsϕ�jJ:�^�ON�YpD��Յ˹?q��B0~�i� ���s{DG�v�7�vU,�=��0������]��VtdD�:��L��̯IG��(DA8\�a&�݋�e�(F|�	��pB#b"�I(��x�ˣݎU節jN�Us-�(�(�{��=ks��������dM�ϻ!�O��ϣ7g��]�l�W�$GV��GH��ګ7��o�߉�3{��k��W�2B�hEx��bw�UGZ��+�F]m܃��&{�[<�p��!A���@�i��LL��ܧ�S��9�^]ΐ�Ia�
c`�0�<��j��܉*�57��y����U�\�
�Q�1؎���N�JV��N�j���R�{K����_��	G��aPDB��
����?O������Z�����wM�P��϶���� (��`�JfDJQQ�Te�������	�JZEiPT�Q���cã"MBD!IT�Д��ۣi�h�r@@�U��T]�W!S�0�E2��0@J�B���0AYXFU dYB!
�P`�B	%��`���JA�e  $�"AG3PkqhUF�Ho�玺������/;�%PDB���6׻�3�n<��.�*ѕ�X;v�T?M`���?�dc���ذ^
B����=LV��"���_ �A���_��"!����C�P�{>'��>��]���É����� ����So���
�"�'��a��mA�g�����c����a���3��m����po��5e����~N�����Tp�V"I$J* %1U
P� %�BJ"R�D�H R 5���*40�3
��D�ECAH� TT�,C@�BHB�P�D�4�)�EhA�% �$�`� aHG�DS !A�`APA�BPA�PA�YARA�BA�YAIA XAe�` Y$AP�i%F�JF ( T
 @h�P�R�(FdDhQ�B�)A�@��&'��A�U�V���bAA��o�����m�|�84�����_������@%I�_����|߁�v���O���{��p��q�� �˱���_����*�g���>_g�������v/�������
���cs���>f����y|C�yx�C����dPDC�Q�7�~�������ߠ}�&�UB��T�?�d��Ooט�'@&w6O��m�l�o��DC}��(�L����?��g�T����Ƌ$�a���g�p��6�?I��u��"�����'��ED?g�|���_���DA<d����������v��=5���y�}���Oן"O����ﰨ"!x)�i��~h����6 A>;�����s���xx>�w?^�	������h�|��8>���.�ߏ�w/�����PDC^}�=v�0��� ��6��G��gӱ�@A0��8ln>�������ePDC�Y?Pǹ��������UD=盰h�	�olx�{�OS~cd�����']�����"�(Hb-n��